
-- Add other necessary VHDL library and use statements here

entity LutROM is
    Port (
        address   : in std_logic_vector(11 downto 0);
        data_out  : out std_logic_vector(1 downto 0)
    );
end LutROM;

architecture Behavioral of LutROM is
    type lut_array is array (natural range <>) of real;
    signal lut : lut_array(0 to 4096 - 1) := ("4.0", "3.6899095998337983", "3.446819498025528", "3.254004476015678", "3.098996239653947", "2.9724968140216057", "2.8675694244650396", "2.7790359972597787", "2.7030285119813557", "2.6366549140818467", "2.577750330836386", "2.524691805726496", "2.4762603299734547", "2.4315380926767896", "2.3898319557366614", "2.3506164566527166", "2.3134913525956295", "2.278149992655911", "2.244355753441236", "2.2119244792824047", "2.1807113940689766", "2.150601343222873", "2.121501515823989", "2.093336013960463", "2.066041798000872", "2.039565656833514", "2.013861941730789", "1.9888908692239768", "1.9646172480600768", "1.9410095223100141", "1.9180390502468643", "1.895679559126896", "1.8739067312818074", "1.852697888305438", "1.8320317485886304", "1.811888239763569", "1.7922483523161437", "1.7730940241229756", "1.7544080482748896", "1.736173998488889", "1.7183761678558405", "1.7009995177475719", "1.6840296345090233", "1.6674526921586128", "1.6512554197652378", "1.6354250725022415", "1.6199494056261248", "1.604816650812377", "1.5900154944185207", "1.5755350573473503", "1.5613648762601824", "1.5474948859474673", "1.5339154027071646", "1.5206171086136226", "1.5075910365840024", "1.4948285561676051", "1.482321359997335", "1.4700614508530614", "1.4580411292946738", "1.4462529818288266", "1.4346898695781471", "1.4233449174254202", "1.4122115036082379", "1.401283249741944", "1.3905540112506531", "1.3800178681876714", "1.3696691164279973", "1.359502259216677", "1.34951199905778", "1.3396932299295938", "1.330041029812404", "1.320550653515895", "1.3112175257938385", "1.3020372347342923", "1.293005525414078", "1.2841182938067772", "1.2753715809339754", "1.2667615672498915", "1.2582845672499712", "1.2499370242943924", "1.2417155056378226", "1.2336166976571104", "1.2256374012689426", "1.2177745275298228", "1.2100250934110284", "1.2023862177415194", "1.1948551173120352", "1.1874291031339104", "1.180105576846386", "1.1728820272664517", "1.1657560270754979", "1.158725229637279", "1.1517873659419173", "1.144940241670891", "1.1381817343781455", "1.131509790782673", "1.1249224241680875", "1.1184177118848995", "1.1119937929513788", "1.1056488657490473", "1.0993811858090086", "1.0931890636854773", "1.0870708629130097", "1.081024998044088", "1.0750499327638299", "1.0691441780787492", "1.06330629057659", "1.057534870754397", "1.0518285614120897", "1.0461860461089187", "1.0406060476802923", "1.0350873268125562", "1.0296286806734123", "1.024228941595751", "1.018886975812767", "1.0136016822423048", "1.0083719913184745", "1.003196863868647", "0.998075290034019", "0.993006288232013", "0.9879889041588388", "0.9830222098306205", "0.9781053026615508", "0.9732373045775984", "0.9684173611643497", "0.9636446408476357", "0.9589183341056257", "0.9542376527111514", "0.9496018290030493", "0.9450101151853738", "0.9404617826533725", "0.9359561213451633", "0.9314924391180897", "0.9270700611487824", "0.9226883293559804", "0.9183466018452162", "0.9140442523744958", "0.9097806698401447", "0.9055552577820225", "0.9013674339073389", "0.8972166296323393", "0.8931022896411536", "0.8890238714611283", "0.8849808450539993", "0.8809726924222725", "0.8769989072302214", "0.8730589944389229", "0.8691524699547791", "0.865278860290999", "0.8614377022415256", "0.8576285425669294", "0.8538509376917889", "0.850104453413117", "0.8463886646193972", "0.8427031550198163", "0.8390475168832945", "0.8354213507869327", "0.8318242653735086", "0.8282558771176691", "0.8247158101004834", "0.821203695792029", "0.8177191728417001", "0.8142618868759413", "0.8108314903031153", "0.8074276421252317", "0.8040500077562717", "0.8006982588468526", "0.7973720731149899", "0.7940711341827217", "0.7907951314183697", "0.7875437597842223", "0.7843167196894294", "0.7811137168479128", "0.7779344621410977", "0.7747786714852845", "0.771646065703481", "0.768536370401528", "0.7654493158483545", "0.7623846368602067", "0.7593420726886994", "0.7563213669125459", "0.7533222673328295", "0.7503445258716814", "0.7473878984742377", "0.7444521450137538", "0.7415370291997563", "0.7386423184891219", "0.7357677839999717", "0.7329132004282772", "0.7300783459670787", "0.7272630022282186", "0.7244669541664971", "0.7216899900061602", "0.7189319011696372", "0.716192482208442", "0.7134715307361625", "0.710768847363459", "0.7080842356350012", "0.705417501968273", "0.7027684555941768", "0.7001369084993734", "0.6975226753702959", "0.6949255735387749", "0.6923454229292231", "0.6897820460073167", "0.687235267730128", "0.6847049154976511", "0.6821908191056777", "0.6796928106999722", "0.6772107247317011", "0.6747443979140748", "0.6722936691801574", "0.6698583796418067", "0.6674383725497037", "0.6650334932544353", "0.6626435891685937", "0.660268509729858", "0.6579081063650267", "0.6555622324549657", "0.653230743300444", "0.6509134960888256", "0.6486103498615923", "0.6463211654826645", "0.6440458056075001", "0.6417841346529415", "0.6395360187677877", "0.6373013258040692", "0.6350799252890016", "0.6328716883975969", "0.6306764879259107", "0.6284941982649067", "0.6263246953749183", "0.6241678567606871", "0.6220235614469631", "0.6198916899546479", "0.6177721242774631", "0.6156647478591293", "0.6135694455710413", "0.6114861036904202", "0.6094146098789334", "0.6073548531617647", "0.605306723907124", "0.6032701138061792", "0.6012449158534052", "0.5992310243273301", "0.597228334771673", "0.5952367439768582", "0.5932561499618986", "0.5912864519566352", "0.5893275503843232", "0.587379346844557", "0.5854417440965214", "0.583514646042564", "0.5815979577120766", "0.579691585245679", "0.5777954358796971", "0.5759094179309274", "0.5740334407816794", "0.5721674148650902", "0.5703112516507024", "0.5684648636303012", "0.5666281643040014", "0.5648010681665785", "0.5629834906940397", "0.5611753483304265", "0.5593765584748446", "0.5575870394687146", "0.5558067105832394", "0.5540354920070818", "0.5522733048342474", "0.5505200710521693", "0.5487757135299881", "0.5470401560070246", "0.5453133230814374", "0.5435951401990665", "0.541885533642453", "0.5401844305200345", "0.5384917587555121", "0.5368074470773827", "0.5351314250086372", "0.5334636228566155", "0.5318039717030205", "0.5301524033940843", "0.528508850530884", "0.5268732464598044", "0.5252455252631446", "0.5236256217498652", "0.5220134714464734", "0.5204090105880427", "0.5188121761093657", "0.5172229056362367", "0.5156411374768604", "0.5140668106133857", "0.5124998646935632", "0.5109402400225203", "0.5093878775546555", "0.5078427188856477", "0.5063047062445782", "0.5047737824861652", "0.5032498910831057", "0.5017329761185256", "0.5002229822785347", "0.4987198548448847", "0.4972235396877288", "0.49573398325848084", "0.4942511325827726", "0.49277493525350624", "0.49130533942400284", "0.4898422938012421", "0.4883857476391946", "0.48693565073224265", "0.4854919534086907", "0.48405460652436083", "0.482623561456275", "0.48119877009642065", "0.47978018484559803", "0.47836775860735015", "0.4769614447819714", "0.4755611972605955", "0.47416697041936007", "0.47277871911364805", "0.47139639867240335", "0.47001996489252085", "0.46864937403330836", "0.46728458281102014", "0.46592554839346195", "0.46457222839466306", "0.463224580869619", "0.46188256430909985", "0.4605461376345251", "0.4592152601929044", "0.45788989175184136", "0.456569992494602", "0.4552555230152442", "0.45394644431380954", "0.4526427177915756", "0.45134430524636765", "0.4500511688679289", "0.4487632712333495", "0.4474805753025522", "0.4462030444138344", "0.4449306422794653", "0.44366333298133936", "0.4424010809666813", "0.4411438510438069", "0.4398916083779342", "0.43864431848704777", "0.4374019472378135", "0.43616446084154414", "0.43493182585021356", "0.4337040091525213", "0.4324809779700044", "0.43126269985319754", "0.4300491426778397", "0.42884027464112773", "0.4276360642580151", "0.42643648035755627", "0.42524149207929557", "0.4240510688696998", "0.42286518047863403", "0.42168379695588126", "0.42050688864770286", "0.4193344261934418", "0.4181663805221665", "0.41700272284935547", "0.415843424673622", "0.4146884577734783", "0.413537794204139", "0.4123914062943625", "0.4112492666433312", "0.410111348117569", "0.40897762384789543", "0.40784806722641687", "0.406722651903554", "0.4056013517851041", "0.4044841410293398", "0.4033709940441415", "0.4022618854841644", "0.40115679024804024", "0.40005568347561127", "0.3989585405451978", "0.3978653370708989", "0.3967760488999242", "0.3956906521099586", "0.3946091230065578", "0.3935314381205747", "0.39245757420561705", "0.39138750823553486", "0.3903212174019377", "0.38925867911174217", "0.38819987098474706", "0.38714477085123916", "0.38609335674962564", "0.3850456069240965", "0.38400149982231235", "0.3829610140931219", "0.3819241285843049", "0.3808908223403427", "0.37986107460021445", "0.37883486479522005", "0.3778121725468285", "0.3767929776645516", "0.3757772601438433", "0.37476500016402253", "0.3737561780862225", "0.3727507744513625", "0.37174876997814466", "0.3707501455610735", "0.36975488226849956", "0.3687629613406858", "0.36777436418789666", "0.3667890723885095", "0.36580706768714866", "0.36482833199284126", "0.3638528473771947", "0.36288059607259554", "0.3619115604704295", "0.36094572311932244", "0.3599830667234021", "0.3590235741405802", "0.3580672283808545", "0.3571140126046308", "0.3561639101210652", "0.3552169043864248", "0.35427297900246846", "0.3533321177148464", "0.3523943044115178", "0.351459523121188", "0.3505277580117632", "0.34959899338882405", "0.3486732136941155", "0.3477504035040568", "0.34683054752826636", "0.34591363060810565", "0.34499963771523917", "0.34408855395021204", "0.3431803645410429", "0.3422750548418346", "0.3413726103314008", "0.3404730166119076", "0.33957625940753244", "0.3386823245631378", "0.3377911980429603", "0.3369028659293156", "0.3360173144213181", "0.33513452983361547", "0.3342544985951379", "0.33337720724786235", "0.33250264244559063", "0.3316307909527421", "0.3307616396431601", "0.3298951754989326", "0.3290313856092263", "0.3281702571691341", "0.327311777478537", "0.32645593394097766", "0.3256027140625479", "0.32475210545079", "0.32390409581360846", "0.32305867295819685", "0.3222158247899756", "0.32137553931154245", "0.3205378046216351", "0.31970260891410635", "0.3188699404769105", "0.31803978769110114", "0.3172121390298423", "0.3163869830574288", "0.31556430842831956", "0.3147441038861813", "0.31392635826294385", "0.31311106047786597", "0.3122981995366118", "0.311487764530339", "0.31067974463479586", "0.30987412910943035", "0.30907090729650877", "0.30827006862024425", "0.30747160258593625", "0.3066754987791189", "0.30588174686472014", "0.30509033658622986", "0.304301257764878", "0.3035145002988221", "0.3027300541623442", "0.3019479094050566", "0.30116805615111775", "0.30039048459845585", "0.2996151850180024", "0.29884214775293444", "0.2980713632179251", "0.2973028218984027", "0.29653651434981937", "0.29577243119692687", "0.2950105631330611", "0.29425090091943573", "0.2934934353844421", "0.29273815742295917", "0.29198505799566987", "0.29123412812838634", "0.2904853589113819", "0.2897387414987318", "0.28899426710766063", "0.2882519270178976", "0.28751171257103914", "0.2867736151699189", "0.28603762627798485", "0.28530373741868337", "0.2845719401748506", "0.283842226188111", "0.283114587158282", "0.28238901484278645", "0.2816655010560706", "0.2809440376690302", "0.2802246166084416", "0.2795072298564008", "0.2787918694497676", "0.27807852747961687", "0.2773671960906961", "0.2766578674808888", "0.2759505339006837", "0.2752451876526513", "0.274541821090925", "0.27384042662068814", "0.27314099669766856", "0.27244352382763665", "0.27174800056591086", "0.27105441951686765", "0.27036277333345793", "0.26967305471672826", "0.26898525641534793", "0.2682993712251414", "0.2676153919886255", "0.2669333115945526", "0.2662531229774587", "0.2655748191172162", "0.2648983930385923", "0.26422383781081255", "0.2635511465471284", "0.2628803124043905", "0.2622113285826268", "0.2615441883246245", "0.26087888491551814", "0.260215411682381", "0.2595537619938221", "0.25889392925958693", "0.25823590693016374", "0.25757968849639273", "0.2569252674890813", "0.2562726374786222", "0.25562179207461744", "0.25497272492550466", "0.2543254297181894", "0.25367990017768033", "0.2530361300667293", "0.25239411318547483", "0.2517538433710902", "0.25111531449743485", "0.25047852047471036", "0.24984345524911972", "0.2492101128025306", "0.24857848715214265", "0.2479485723501581", "0.24732036248345635", "0.24669385167327187", "0.24606903407487613", "0.24544590387726287", "0.24482445530283664", "0.24420468260710515", "0.24358658007837503", "0.24297014203745074", "0.242355362837337", "0.2417422368629444", "0.24113075853079877", "0.24052092228875294", "0.23991272261570207", "0.2393061540213028", "0.2387012110456944", "0.2380978882592238", "0.23749618026217323", "0.23689608168449117", "0.23629758718552613", "0.23570069145376332", "0.23510538920656446", "0.23451167518991", "0.23391954417814498", "0.2333289909737267", "0.232740010406976", "0.2321525973358307", "0.23156674664560242", "0.23098245324873512", "0.23039971208456717", "0.2298185181190958", "0.2292388663447434", "0.22866075178012799", "0.2280841694698343", "0.22750911448418898", "0.22693558191903707", "0.22636356689552176", "0.225793064559866", "0.22522407008315676", "0.22465657866113187", "0.22409058551396838", "0.22352608588607417", "0.2229630750458814", "0.22240154828564196", "0.22184150092122562", "0.22128292829192003", "0.22072582576023328", "0.22017018871169805", "0.21961601255467825", "0.2190632927201776", "0.21851202466165065", "0.2179622038548154", "0.21741382579746793", "0.21686688600929935", "0.21632138003171453", "0.21577730342765303", "0.21523465178141143", "0.21469342069846797", "0.21415360580530934", "0.21361520274925846", "0.2130782071983051", "0.2125426148409374", "0.21200842138597625", "0.21147562256241031", "0.21094421411923348", "0.21041419182528429", "0.20988555146908583", "0.20935828885868932", "0.20883239982151744", "0.20830788020421037", "0.20778472587247346", "0.20726293271092594", "0.2067424966229518", "0.20622341353055199", "0.20570567937419834", "0.20518929011268872", "0.20467424172300405", "0.20416053020016678", "0.2036481515571007", "0.20313710182449232", "0.20262737705065367", "0.20211897330138678", "0.20161188665984914", "0.20110611322642089", "0.2006016491185734", "0.20009849047073905", "0.19959663343418277", "0.1990960741768742", "0.1985968088833619", "0.19809883375464854", "0.1976021450080674", "0.19710673887716024", "0.19661261161155635", "0.1961197594768531", "0.19562817875449712", "0.19513786574166753", "0.19464881675115978", "0.19416102811127098", "0.1936744961656862", "0.1931892172733661", "0.1927051878084358", "0.19222240416007458", "0.191740862732407", "0.19126055994439517", "0.19078149222973173", "0.19030365603673435", "0.18982704782824128", "0.18935166408150758", "0.18887750128810282", "0.18840455595380967", "0.18793282459852348", "0.187462303756153", "0.18699298997452177", "0.1865248798152713", "0.18605796985376416", "0.18559225667898888", "0.18512773689346548", "0.18466440711315193", "0.18420226396735176", "0.18374130409862213", "0.18328152416268362", "0.1828229208283301", "0.18236549077734007", "0.18190923070438844", "0.18145413731695959", "0.18100020733526123", "0.1805474374921388", "0.180095824532991", "0.1796453652156862", "0.17919605631047955", "0.17874789459993082", "0.1783008768788233", "0.17785499995408338", "0.1774102606447008", "0.17696665578164994", "0.1765241822078116", "0.1760828367778959", "0.1756426163583655", "0.17520351782735988", "0.17476553807462036", "0.17432867400141566", "0.17389292252046842", "0.17345828055588222", "0.17302474504306928", "0.17259231292867927", "0.1721609811705283", "0.17173074673752883", "0.17130160660962032", "0.17087355777770044", "0.1704465972435569", "0.17002072201980006", "0.16959592912979624", "0.16917221560760123", "0.16874957849789518", "0.16832801485591734", "0.16790752174740184", "0.16748809624851435", "0.16706973544578846", "0.16665243643606362", "0.16623619632642297", "0.1658210122341324", "0.1654068812865794", "0.1649938006212131", "0.16458176738548475", "0.1641707787367886", "0.16376083184240334", "0.16335192387943429", "0.162944052034756", "0.1625372135049553", "0.162131405496275", "0.16172662522455794", "0.16132286991519212", "0.16092013680305534", "0.16051842313246129", "0.16011772615710565", "0.15971804314001273", "0.15931937135348295", "0.15892170807904002", "0.1585250506073795", "0.15812939623831734", "0.15773474228073883", "0.1573410860525483", "0.15694842488061894", "0.1565567561007436", "0.15616607705758534", "0.1557763851046289", "0.1553876776041325", "0.15499995192708016", "0.15461320545313406", "0.1542274355705879", "0.15384263967632014", "0.15345881517574794", "0.15307595948278174", "0.15269407001977958", "0.15231314421750222", "0.1519331795150691", "0.15155417335991359", "0.15117612320773968", "0.15079902652247854", "0.15042288077624555", "0.15004768344929764", "0.1496734320299911", "0.14930012401473974", "0.1489277569079735", "0.14855632822209702", "0.1481858354774491", "0.1478162762022623", "0.14744764793262247", "0.1470799482124296", "0.14671317459335784", "0.14634732463481667", "0.1459823959039124", "0.14561838597540921", "0.14525529243169147", "0.14489311286272583", "0.14453184486602383", "0.1441714860466046", "0.14381203401695822", "0.1434534863970091", "0.14309584081407978", "0.14273909490285488", "0.1423832463053457", "0.14202829267085484", "0.14167423165594092", "0.1413210609243842", "0.14096877814715172", "0.14061738100236343", "0.1402668671752582", "0.13991723435816006", "0.13956848025044497", "0.13922060255850768", "0.1388735989957289", "0.13852746728244278", "0.1381822051459045", "0.1378378103202585", "0.13749428054650623", "0.13715161357247516", "0.13680980715278693", "0.13646885904882694", "0.13612876702871296", "0.13578952886726497", "0.13545114234597472", "0.13511360525297564", "0.13477691538301295", "0.13444107053741433", "0.13410606852406007", "0.13377190715735449", "0.13343858425819646", "0.13310609765395107", "0.1327744451784211", "0.1324436246718185", "0.1321136339807367", "0.13178447095812254", "0.1314561334632487", "0.13112861936168627", "0.1308019265252777", "0.13047605283210942", "0.1301509961664855", "0.12982675441890065", "0.12950332548601415", "0.1291807072706233", "0.12885889768163783", "0.12853789463405355", "0.1282176960489272", "0.12789829985335083", "0.12757970398042634", "0.12726190636924073", "0.12694490496484112", "0.1266286977182098", "0.12631328258624008", "0.12599865753171158", "0.1256848205232663", "0.12537176953538456", "0.12505950254836104", "0.12474801754828121", "0.124437312526998", "0.12412738548210799", "0.12381823441692882", "0.1235098573404757", "0.12320225226743903", "0.12289541721816118", "0.12258935021861449", "0.12228404930037848", "0.12197951250061793", "0.12167573786206078", "0.12137272343297589", "0.12107046726715179", "0.12076896742387476", "0.12046822196790727", "0.12016822896946702", "0.11986898650420551", "0.11957049265318691", "0.1192727455028676", "0.11897574314507485", "0.11867948367698672", "0.11838396520111132", "0.11808918582526648", "0.11779514366255951", "0.11750183683136742", "0.11720926345531664", "0.11691742166326333", "0.11662630958927372", "0.11633592537260473", "0.11604626715768403", "0.11575733309409143", "0.11546912133653911", "0.11518163004485293", "0.11489485738395347", "0.1146088015238369", "0.11432346063955677", "0.11403883291120516", "0.11375491652389412", "0.11347170966773767", "0.11318921053783328", "0.11290741733424382", "0.11262632826197978", "0.1123459415309812", "0.11206625535609971", "0.1117872679570813", "0.11150897755854851", "0.11123138238998288", "0.11095448068570789", "0.11067827068487154", "0.11040275063142913", "0.11012791877412653", "0.10985377336648304", "0.10958031266677447", "0.10930753493801675", "0.10903543844794893", "0.10876402146901694", "0.10849328227835711", "0.10822321915777965", "0.10795383039375252", "0.1076851142773855", "0.10741706910441391", "0.10714969317518254", "0.10688298479463021", "0.10661694227227354", "0.1063515639221916", "0.10608684806301026", "0.10582279301788643", "0.10555939711449307", "0.10529665868500357", "0.10503457606607654", "0.10477314759884078", "0.10451237162888022", "0.10425224650621866", "0.10399277058530526", "0.10373394222499957", "0.1034757597885565", "0.1032182216436122", "0.10296132616216923", "0.10270507172058187", "0.10244945669954203", "0.10219447948406483", "0.10194013846347416", "0.10168643203138873", "0.10143335858570794", "0.10118091652859759", "0.10092910426647635", "0.10067792021000144", "0.10042736277405521", "0.10017743037773123", "0.09992812144432049", "0.0996794344012981", "0.09943136768030965", "0.09918391971715765", "0.09893708895178828", "0.09869087382827807", "0.09844527279482071", "0.09820028430371369", "0.09795590681134544", "0.09771213877818208", "0.09746897866875459", "0.09722642495164595", "0.09698447609947802", "0.0967431305888991", "0.09650238690057114", "0.09626224351915684", "0.09602269893330738", "0.09578375163564985", "0.09554540012277453", "0.09530764289522284", "0.09507047845747488", "0.09483390531793687", "0.09459792198892941", "0.09436252698667513", "0.09412771883128634", "0.0938934960467534", "0.09365985716093254", "0.0934268007055338", "0.09319432521610944", "0.09296242923204201", "0.09273111129653243", "0.09250036995658864", "0.09227020376301359", "0.09204061127039394", "0.09181159103708841", "0.09158314162521616", "0.09135526160064565", "0.09112794953298312", "0.09090120399556113", "0.09067502356542749", "0.090449406823334", "0.09022435235372533", "0.08999985874472764", "0.08977592458813795", "0.08955254847941264", "0.08932972901765693", "0.08910746480561371", "0.08888575444965263", "0.08866459655975953", "0.08844398974952546", "0.08822393263613593", "0.08800442384036046", "0.08778546198654179", "0.08756704570258522", "0.08734917361994836", "0.08713184437363028", "0.08691505660216134", "0.0866988089475927", "0.08648310005548603", "0.086267928574903", "0.08605329315839524", "0.08583919246199415", "0.08562562514520038", "0.08541258987097411", "0.08520008530572477", "0.08498811011930091", "0.08477666298498039", "0.08456574257946024", "0.0843553475828469", "0.08414547667864625", "0.08393612855375368", "0.08372730189844453", "0.08351899540636415", "0.0833112077745182", "0.083103937703263", "0.08289718389629598", "0.08269094506064599", "0.08248521990666365", "0.08228000714801206", "0.0820753055016571", "0.0818711136878582", "0.08166743043015874", "0.08146425445537671", "0.08126158449359557", "0.08105941927815476", "0.08085775754564045", "0.08065659803587645", "0.080455939491915", "0.08025578066002743", "0.0800561202896954", "0.07985695713360144", "0.0796582899476203", "0.07946011749080951", "0.07926243852540092", "0.07906525181679128", "0.07886855613353365", "0.07867235024732849", "0.07847663293301471", "0.07828140296856095", "0.07808665913505691", "0.07789240021670439", "0.07769862500080887", "0.07750533227777057", "0.07731252084107605", "0.07712018948728956", "0.07692833701604428", "0.07673696223003405", "0.07654606393500482", "0.07635564093974596", "0.07616569205608202", "0.07597621609886443", "0.07578721188596275", "0.07559867823825675", "0.07541061397962781", "0.07522301793695069", "0.07503588894008534", "0.07484922582186872", "0.07466302741810636", "0.07447729256756455", "0.07429202011196194", "0.07410720889596147", "0.07392285776716243", "0.07373896557609232", "0.07355553117619872", "0.0733725534238416", "0.07319003117828499", "0.07300796330168938", "0.07282634865910359", "0.07264518611845704", "0.07246447455055172", "0.07228421282905459", "0.07210439983048969", "0.07192503443423025", "0.0717461155224912", "0.07156764198032117", "0.0713896126955951", "0.07121202655900641", "0.0710348824640593", "0.07085817930706133", "0.07068191598711575", "0.07050609140611387", "0.07033070446872772", "0.07015575408240239", "0.06998123915734854", "0.0698071586065351", "0.06963351134568171", "0.06946029629325133", "0.06928751237044296", "0.06911515850118426", "0.06894323361212407", "0.06877173663262534", "0.06860066649475773", "0.0684300221332903", "0.0682598024856844", "0.0680900064920865", "0.06792063309532079", "0.06775168124088224", "0.0675831498769294", "0.06741503795427725", "0.06724734442639019", "0.06708006824937486", "0.06691320838197327", "0.0667467637855556", "0.06658073342411337", "0.06641511626425232", "0.0662499112751856", "0.06608511742872683", "0.06592073369928299", "0.06575675906384784", "0.06559319250199488", "0.06543003299587051", "0.06526727953018738", "0.06510493109221732", "0.06494298667178487", "0.06478144526126033", "0.06462030585555303", "0.06445956745210482", "0.06429922905088319", "0.06413928965437458", "0.063979748267578", "0.06382060389799811", "0.06366185555563875", "0.06350350225299638", "0.06334554300505359", "0.06318797682927225", "0.06303080274558741", "0.06287401977640053", "0.06271762694657305", "0.06256162328341999", "0.0624060078167035", "0.06225077957862635", "0.062095937603825695", "0.06194148092936652", "0.06178740859473548", "0.061633719641834325", "0.06148041311497384", "0.06132748806086726", "0.06117494352862436", "0.06102277856974477", "0.06087099223811209", "0.060719583589987414", "0.06056855168400332", "0.06041789558115748", "0.060267614344806854", "0.06011770704066095", "0.05996817273677639", "0.059819010503550256", "0.05967021941371422", "0.05952179854232852", "0.05937374696677576", "0.05922606376675503", "0.05907874802427567", "0.05893179882365163", "0.05878521525149501", "0.05863899639671054", "0.0584931413504893", "0.05834764920630306", "0.058202519059898115", "0.058057750009289616", "0.0579133411547555", "0.057769291598830846", "0.05762560044630177", "0.05748226680419987", "0.057339289781796185", "0.057196668490595515", "0.05705440204433073", "0.056912489558956815", "0.05677093015264534", "0.0566297229457785", "0.056488867060943734", "0.05634836162292766", "0.056208205758710716", "0.05606839859746129", "0.055928939270530234", "0.055789826911445066", "0.05565106065590465", "0.05551263964177324", "0.055374563009075194", "0.05523682989998925", "0.0550994394588431", "0.054962390832107744", "0.0548256831683921", "0.054689315618437415", "0.05455328733511177", "0.05441759747340482", "0.05428224519042203", "0.05414722964537951", "0.05401254999959841", "0.0538782054164997", "0.053744195061598575", "0.05361051810249932", "0.053477173708889665", "0.05334416105253582", "0.05321147930727676", "0.053079127649019196", "0.0529471052557321", "0.05281541130744162", "0.05268404498622554", "0.05255300547620837", "0.052422291963555814", "0.05229190363646961", "0.05216183968518256", "0.05203209930195299", "0.05190268168105986", "0.05177358601879737", "0.05164481151347004", "0.051516357365387344", "0.05138822277685885", "0.05126040695218885", "0.05113290909767146", "0.05100572842158543", "0.05087886413418919", "0.05075231544771567", "0.05062608157636742", "0.05050016173631141", "0.050374555145674245", "0.05024926102453694", "0.05012427859493007", "0.049999607080828845", "0.04987524570814803", "0.04975119370473715", "0.049627450300375374", "0.04950401472676692", "0.04938088621753573", "0.04925806400822104", "0.049135547336272116", "0.04901333544104371", "0.04889142756379095", "0.04876982294766478", "0.04864852083770685", "0.04852752048084503", "0.048406821125888316", "0.0482864220235223", "0.0481663224263042", "0.04804652158865831", "0.04792701876687109", "0.047807813219086503", "0.0476889042053014", "0.0475702909873606", "0.04745197282895248", "0.047333948995604024", "0.04721621875467641", "0.047098781375360145", "0.046981636128670595", "0.04686478228744324", "0.04674821912632924", "0.04663194592179049", "0.04651596195209553", "0.04640026649731449", "0.046284858839314866", "0.046169738261756736", "0.04605490405008844", "0.045940355491541886", "0.04582609187512805", "0.04571211249163267", "0.04559841663361147", "0.04548500359538592", "0.04537187267303858", "0.04525902316440884", "0.04514645436908833", "0.04503416558841659", "0.04492215612547651", "0.044810425285090175", "0.044698972373814205", "0.044587796699935546", "0.044476897573467004", "0.044366274306142976", "0.04425592621141498", "0.04414585260444754", "0.044036052802113555", "0.0439265261229902", "0.04381727188735468", "0.043708289417179684", "0.0435995780361294", "0.04349113706955498", "0.043382965844490536", "0.04327506368964865", "0.04316742993541644", "0.043060063913850984", "0.042952964958675434", "0.042846132405274566", "0.04273956559069081", "0.042633263853619846", "0.042527226534406694", "0.042421452975041275", "0.0423159425191546", "0.04221069451201426", "0.04210570830052065", "0.042000983233202616", "0.041896518660213454", "0.041792313933326886", "0.0416883684059328", "0.04158468143303338", "0.04148125237123888", "0.04137808057876376", "0.04127516541542243", "0.04117250624262543", "0.041070102423375256", "0.040967953322262496", "0.04086605830546168", "0.04076441674072749", "0.040663027997390584", "0.04056189144635379", "0.040461006460088045", "0.04036037241262856", "0.04025998867957078", "0.040159854638066504", "0.04005996966682006", "0.03996033314608421", "0.03986094445765651", "0.03976180298487519", "0.039662908112615455", "0.03956425922728549", "0.03946585571682277", "0.039367696970690036", "0.03926978237987163", "0.03917211133686954", "0.03907468323569974", "0.0389774974718882", "0.03888055344246728", "0.0387838505459718", "0.038687388182435396", "0.03859116575338664", "0.038495182661845366", "0.038399438312318984", "0.03830393211079851", "0.03820866346475519", "0.03811363178313647", "0.038018836476362505", "0.03792427695632233", "0.03782995263637029", "0.03773586293132223", "0.03764200725745204", "0.037548385032487724", "0.03745499567560801", "0.03736183860743852", "0.037268913250048295", "0.03717621902694604", "0.03708375536307665", "0.03699152168481746", "0.03689951741997486", "0.036807741997780495", "0.036716194848887794", "0.03662487540536846", "0.036533783100708817", "0.036442917369806344", "0.03635227764896604", "0.0362618633758971", "0.036171673989709094", "0.03608170893090878", "0.03599196764139635", "0.03590244956446212", "0.035813154144782894", "0.035724080828418665", "0.03563522906280894", "0.03554659829676957", "0.035458187980488984", "0.03536999756552501", "0.03528202650480129", "0.03519427425260392", "0.03510674026457811", "0.0350194239977246", "0.03493232491039648", "0.034845442462295616", "0.03475877611446947", "0.034672325329307516", "0.034586089570538076", "0.03450006830322483", "0.03441426099376359", "0.034328667109878815", "0.03424328612062054", "0.03415811749636074", "0.0340731607087903", "0.03398841523091554", "0.03390388053705504", "0.033819556102836254", "0.03373544140519232", "0.03365153592235878", "0.03356783913387027", "0.033484350520557364", "0.03340106956454323", "0.0333179957492405", "0.033235128559347925", "0.03315246748084732", "0.03307001200100019", "0.03298776160834468", "0.03290571579269221", "0.03282387404512456", "0.03274223585799037", "0.032660800724902225", "0.03257956814073338", "0.03249853760161465", "0.03241770860493123", "0.03233708064931962", "0.032256653234664485", "0.03217642586209538", "0.032096398033983974", "0.03201656925394059", "0.03193693902681138", "0.03185750685867502", "0.03177827225683985", "0.03169923472984058", "0.03162039378743547", "0.03154174894060301", "0.0314632997015391", "0.03138504558365385", "0.03130698610156868", "0.031229120771113145", "0.031151449109322084", "0.031073970634432447", "0.030996684865880468", "0.030919591324298494", "0.0308426895315121", "0.030765979010537133", "0.03068945928557663", "0.030613129882018", "0.030536990326429893", "0.03046104014655948", "0.03038527887132923", "0.030309706030834254", "0.030234321156339165", "0.0301591237802753", "0.030084113436237694", "0.030009289658982297", "0.02993465198442294", "0.029860199949628616", "0.029785933092820398", "0.029711850953368747", "0.029637953071790506", "0.029564238989746115", "0.029490708250036756", "0.029417360396601453", "0.02934419497451432", "0.02927121152998161", "0.029198409610339038", "0.02912578876404882", "0.029053348540696963", "0.028981088490990393", "0.028909008166754232", "0.0288371071209289", "0.02876538490756752", "0.028693841081832858", "0.028622475199994876", "0.02855128681942771", "0.02848027549860708", "0.028409440797107426", "0.02833878227559929", "0.028268299495846465", "0.028197992020703312", "0.028127859414112125", "0.028057901241100247", "0.02798811706777753", "0.02791850646133351", "0.027849068990034805", "0.027779804223222366", "0.027710711731308856", "0.027641791085775892", "0.027573041859171518", "0.027504463625107375", "0.027436055958256204", "0.027367818434349076", "0.027299750630172856", "0.027231852123567477", "0.02716412249342344", "0.02709656131967903", "0.02702916818331782", "0.026961942666366076", "0.026894884351890063", "0.026827992823993556", "0.026761267667815156", "0.026694708469525808", "0.026628314816326118", "0.026562086296443937", "0.026496022499131622", "0.026430123014663638", "0.026364387434333895", "0.026298815350453298", "0.02623340635634713", "0.026168160046352612", "0.02610307601581627", "0.026038153861091578", "0.025973393179536265", "0.025908793569509928", "0.025844354630371536", "0.025780075962476865", "0.02571595716717612", "0.025651997846811336", "0.02558819760471402", "0.02552455604520258", "0.025461072773580003", "0.025397747396131223", "0.02533457952012085", "0.02527156875379058", "0.025208714706356893", "0.025146016988008495", "0.02508347520990404", "0.02502108898416956", "0.024958857923896183", "0.02489678164313763", "0.02483485975690791", "0.024773091881178846", "0.024711477632877718", "0.02465001662988492", "0.024588708491031504", "0.024527552836096932", "0.02446654928580657", "0.02440569746182945", "0.024344996986775835", "0.024284447484194963", "0.02422404857857259", "0.0241637998953288", "0.02410370106081552", "0.024043751702314375", "0.023983951448034193", "0.023924299927108837", "0.023864796769594805", "0.023805441606469007", "0.023746234069626414", "0.023687173791877774", "0.02362826040694744", "0.02356949354947088", "0.023510872854992648", "0.023452397959963928", "0.023394068501740407", "0.02333588411857992", "0.023277844449640307", "0.02321994913497705", "0.023162197815541193", "0.02310459013317694", "0.023047125730619566", "0.022989804251493114", "0.022932625340308245", "0.022875588642459966", "0.0228186938042255", "0.022761940472762015", "0.02270532829610446", "0.022648856923163454", "0.022592526003722958", "0.02253633518843824", "0.022480284128833593", "0.022424372477300288", "0.022368599887094276", "0.02231296601233421", "0.022257470507999075", "0.022202113029926286", "0.022146893234809346", "0.022091810780195863", "0.022036865324485313", "0.021982056526927005", "0.021927384047617893", "0.021872847547500556", "0.02181844668836098", "0.021764181132826535", "0.021710050544363875", "0.02165605458727681", "0.021602192926704282", "0.021548465228618197", "0.021494871159821464", "0.0214414103879458", "0.021388082581449815", "0.021334887409616792", "0.021281824542552768", "0.021228893651184393", "0.021176094407256964", "0.02112342648333229", "0.021070889552786812", "0.021018483289809365", "0.020966207369399373", "0.020914061467364665", "0.02086204526031957", "0.020810158425682828", "0.020758400641675636", "0.020706771587319674", "0.020655270942435026", "0.020603898387638306", "0.020552653604340554", "0.02050153627474537", "0.02045054608184685", "0.0203996827094277", "0.020348945842057185", "0.020298335165089262", "0.02024785036466055", "0.02019749112768845", "0.020147257141869126", "0.020097148095675647", "0.020047163678355972", "0.019997303579931108", "0.019947567491193106", "0.019897955103703176", "0.019848466109789808", "0.019799100202546778", "0.019749857075831354", "0.01970073642426227", "0.019651737943217954", "0.019602861328834525", "0.019554106278004", "0.019505472488372342", "0.01945695965833766", "0.01940856748704825", "0.019360295674400795", "0.019312143921038447", "0.01926411192834904", "0.01921619939846316", "0.019168406034252374", "0.019120731539327303", "0.019073175618035825", "0.019025737975461296", "0.018978418317420594", "0.018931216350462417", "0.01888413178186536", "0.018837164319636193", "0.01879031367250796", "0.018743579549938244", "0.018696961662107308", "0.018650459719916367", "0.018604073434985692", "0.018557802519652927", "0.01851164668697121", "0.018465605650707477", "0.018419679125340604", "0.018373866826059734", "0.018328168468762396", "0.018282583770052853", "0.018237112447240217", "0.018191754218336825", "0.018146508802056423", "0.018101375917812416", "0.018056355285716162", "0.018011446626575164", "0.017966649661891432", "0.017921964113859698", "0.01787738970536572", "0.01783292615998448", "0.017788573201978644", "0.01774433055629664", "0.017700197948571104", "0.017656175105117123", "0.017612261752930552", "0.017568457619686246", "0.017524762433736546", "0.017481175924109384", "0.017437697820506703", "0.01739432785330286", "0.01735106575354277", "0.0173079112529404", "0.017264864083877007", "0.017221923979399548", "0.017179090673218912", "0.017136363899708455", "0.017093743393902135", "0.017051228891493023", "0.01700882012883161", "0.016966516842924176", "0.016924318771431128", "0.01688222565266543", "0.016840237225590943", "0.016798353229820817", "0.01675657340561587", "0.016714897493882948", "0.01667332523617339", "0.016631856374681363", "0.01659049065224229", "0.016549227812331205", "0.016508067599061288", "0.016467009757182093", "0.016426054032078138", "0.016385200169767206", "0.016344447916898857", "0.016303797020752755", "0.016263247229237204", "0.016222798290887526", "0.016182449954864512", "0.016142201970952872", "0.01610205408955969", "0.016062006061712812", "0.016022057639059412", "0.01598220857386438", "0.01594245861900876", "0.015902807527988293", "0.015863255054911846", "0.015823800954499874", "0.01578444498208293", "0.015745186893600133", "0.01570602644559762", "0.0156669633952271", "0.015627997500244312", "0.01558912851900754", "0.015550356210476035", "0.015511680334208687", "0.015473100650362335", "0.01543461691969043", "0.015396228903541481", "0.015357936363857606", "0.015319739063172995", "0.015281636764612524", "0.015243629231890229", "0.015205716229307853", "0.015167897521753399", "0.015130172874699612", "0.015092542054202619", "0.015055004826900406", "0.015017560960011413", "0.01498021022133301", "0.014942952379240213", "0.014905787202684057", "0.01486871446119031", "0.014831733924857975", "0.01479484536435789", "0.014758048550931248", "0.014721343256388308", "0.01468472925310682", "0.014648206314030692", "0.014611774212668651", "0.014575432723092677", "0.01453918161993674", "0.014503020678395344", "0.014466949674222145", "0.01443096838372851", "0.014395076583782262", "0.014359274051806124", "0.014323560565776466", "0.014287935904221881", "0.014252399846221824", "0.014216952171405192", "0.014181592659949043", "0.014146321092577168", "0.014111137250558755", "0.014076040915707029", "0.014041031870377902", "0.014006109897468587", "0.013971274780416324", "0.013936526303196986", "0.013901864250323718", "0.013867288406845665", "0.013832798558346597", "0.013798394490943578", "0.013764075991285655", "0.01372984284655254", "0.013695694844453241", "0.013661631773224813", "0.013627653421631004", "0.013593759578960961", "0.013559950035027907", "0.013526224580167867", "0.0134925830052383", "0.013459025101616895", "0.01342555066120023", "0.01339215947640244", "0.013358851340154014", "0.013325626045900454", "0.013292483387601006", "0.013259423159727389", "0.013226445157262522", "0.013193549175699216", "0.013160735011038968", "0.013128002459790651", "0.013095351318969273", "0.013062781386094667", "0.013030292459190358", "0.012997884336782147", "0.01296555681789699", "0.012933309702061692", "0.012901142789301694", "0.012869055880139774", "0.012837048775594894", "0.012805121277180913", "0.01277327318690533", "0.012741504307268165", "0.012709814441260585", "0.012678203392363805", "0.01264667096454781", "0.01261521696227016", "0.012583841190474726", "0.012552543454590604", "0.012521323560530742", "0.012490181314690877", "0.012459116523948256", "0.01242812899566048", "0.01239721853766425", "0.01236638495827426", "0.012335628066281938", "0.012304947670954296", "0.012274343582032743", "0.012243815609731866", "0.012213363564738322", "0.012182987258209611", "0.012152686501772932", "0.012122461107523968", "0.012092310888025825", "0.012062235656307726", "0.01203223522586397", "0.012002309410652726", "0.011972458025094885", "0.011942680884072887", "0.01191297780292962", "0.01188334859746724", "0.011853793083946042", "0.01182431107908331", "0.011794902400052204", "0.01176556686448057", "0.011736304290449886", "0.01170711449649409", "0.011677997301598434", "0.011648952525198413", "0.011619979987178612", "0.011591079507871598", "0.0115622509080568", "0.011533494008959417", "0.011504808632249256", "0.011476194600039704", "0.011447651734886566", "0.011419179859786997", "0.011390778798178349", "0.011362448373937191", "0.011334188411378067", "0.011305998735252527", "0.011277879170747991", "0.011249829543486647", "0.011221849679524415", "0.011193939405349837", "0.01116609854788301", "0.011138326934474512", "0.011110624392904337", "0.011082990751380799", "0.011055425838539508", "0.011027929483442285", "0.01100050151557611", "0.010973141764852026", "0.010945850061604175", "0.01091862623658863", "0.010891470120982438", "0.010864381546382525", "0.01083736034480468", "0.010810406348682458", "0.010783519390866246", "0.010756699304622105", "0.010729945923630791", "0.010703259081986783", "0.010676638614197131", "0.010650084355180528", "0.010623596140266247", "0.01059717380519313", "0.010570817186108535", "0.010544526119567405", "0.010518300442531141", "0.010492139992366681", "0.010466044606845457", "0.010440014124142388", "0.010414048382834865", "0.010388147221901782", "0.010362310480722517", "0.010336537999075933", "0.010310829617139403", "0.010285185175487776", "0.010259604515092446", "0.010234087477320328", "0.010208633903932897", "0.010183243637085159", "0.010157916519324742", "0.010132652393590869", "0.0101074511032134", "0.010082312491911863", "0.010057236403794485", "0.010032222683357203", "0.010007271175482732", "0.009982381725439596", "0.009957554178881148", "0.009932788381844634", "0.009908084180750235", "0.009883441422400089", "0.00985885995397738", "0.009834339623045384", "0.009809880277546475", "0.00978548176580125", "0.009761143936507548", "0.009736866638739522", "0.009712649721946697", "0.009688493035953054", "0.009664396430956065", "0.009640359757525798", "0.009616382866603983", "0.00959246560950308", "0.009568607837905325", "0.009544809403861912", "0.00952107015979194", "0.0094973899584816", "0.009473768653083222", "0.009450206097114375", "0.009426702144456931", "0.009403256649356201", "0.009379869466420011", "0.009356540450617788", "0.009333269457279691", "0.00931005634209567", "0.00928690096111462", "0.009263803170743453", "0.009240762827746232", "0.009217779789243239", "0.009194853912710176", "0.009171985055977163", "0.009149173077227958", "0.00912641783499903", "0.009103719188178691", "0.009081076996006196", "0.009058491118070944", "0.00903596141431151", "0.00901348774501483", "0.008991069970815365", "0.00896870795269415", "0.008946401551978017", "0.008924150630338685", "0.008901955049791925", "0.00887981467269667", "0.008857729361754241", "0.00883569898000738", "0.008813723390839504", "0.008791802457973803", "0.008769936045472415", "0.008748124017735559", "0.008726366239500726", "0.00870466257584183", "0.00868301289216835", "0.008661417054224537", "0.008639874928088521", "0.008618386380171547", "0.008596951277217104", "0.008575569486300118", "0.008554240874826098", "0.008532965310530357", "0.008511742661477164", "0.008490572796058932", "0.008469455582995403", "0.008448390891332837", "0.008427378590443178", "0.00840641855002328", "0.008385510640094074", "0.008364654730999769", "0.008343850693407049", "0.008323098398304274", "0.008302397717000656", "0.008281748521125502", "0.008261150682627392", "0.008240604073773373", "0.008220108567148197", "0.008199664035653522", "0.008179270352507107", "0.00815892739124204", "0.008138635025705963", "0.00811839313006025", "0.008098201578779282", "0.008078060246649628", "0.008057969008769292", "0.0080379277405469", "0.008017936317701", "0.007997994616259205", "0.007978102512557483", "0.00795825988323938", "0.007938466605255238", "0.007918722555861435", "0.007899027612619644", "0.007879381653396062", "0.007859784556360624", "0.007840236199986321", "0.007820736463048353", "0.007801285224623452", "0.007781882364089092", "0.0077625277611227655", "0.007743221295701195", "0.007723962848099667", "0.007704752298891194", "0.007685589528945846", "0.00766647441942998", "0.00764740685180552", "0.007628386707829186", "0.00760941386955181", "0.007590488219317581", "0.007571609639763285", "0.007552778013817659", "0.007533993224700564", "0.007515255155922336", "0.007496563691283033", "0.007477918714871724", "0.007459320111065742", "0.007440767764530033", "0.007422261560216354", "0.007403801383362628", "0.0073853871194922045", "0.007367018654413157", "0.007348695874217553", "0.0073304186652807845", "0.007312186914260837", "0.007294000508097595", "0.007275859334012139", "0.007257763279506054", "0.007239712232360707", "0.0072217060806365856", "0.007203744712672587", "0.007185828017085311", "0.007167955882768396", "0.0071501281988918175", "0.007132344854901199", "0.00711460574051713", "0.007096910745734483", "0.007079259760821716", "0.0070616526763202184", "0.007044089383043618", "0.007026569772077107", "0.007009093734776741", "0.006991661162768833", "0.00697427194794919", "0.006956925982482518", "0.006939623158801726", "0.006922363369607233", "0.006905146507866352", "0.006887972466812595", "0.006870841139945013", "0.006853752421027544", "0.006836706204088355", "0.006819702383419163", "0.006802740853574614", "0.006785821509371605", "0.0067689442458886435", "0.006752108958465172", "0.0067353155427009774", "0.0067185638944554605", "0.0067018539098470655", "0.006685185485252591", "0.006668558517306575", "0.0066519729029006144", "0.0066354285391827745", "0.006618925323556926", "0.006602463153682089", "0.006586041927471859", "0.006569661543093694", "0.006553321898968349", "0.006537022893769216", "0.006520764426421703", "0.006504546396102583", "0.006488368702239431", "0.006472231244509924", "0.006456133922841269", "0.006440076637409571", "0.006424059288639212", "0.006408081777202216", "0.006392144004017669", "0.006376245870251078", "0.006360387277313764", "0.006344568126862261", "0.006328788320797678", "0.006313047761265126", "0.006297346350653092", "0.006281683991592839", "0.006266060586957785", "0.006250476039862933", "0.006234930253664244", "0.006219423131958048", "0.006203954578580447", "0.006188524497606718", "0.0061731327933507016", "0.006157779370364239", "0.00614246413343656", "0.006127186987593696", "0.006111947838097892", "0.006096746590447024", "0.006081583150373996", "0.006066457423846177", "0.006051369317064814", "0.006036318736464424", "0.0060213055887122545", "0.0060063297807076785", "0.005991391219581622", "0.00597648981269599", "0.005961625467643095", "0.005946798092245069", "0.005932007594553314", "0.00591725388284792", "0.005902536865637099", "0.005887856451656597", "0.005873212549869184", "0.005858605069464015", "0.005844033919856124", "0.005829499010685844", "0.005815000251818229", "0.005800537553342528", "0.005786110825571603", "0.005771719979041388", "0.0057573649245103034", "0.005743045572958765", "0.005728761835588555", "0.005714513623822329", "0.005700300849303043", "0.0056861234238934156", "0.005671981259675351", "0.0056578742689494576", "0.0056438023642344255", "0.0056297654582665455", "0.0056157634639991405", "0.005601796294602034", "0.005587863863460993", "0.005573966084177224", "0.005560102870566817", "0.005546274136660194", "0.005532479796701631", "0.005518719765148653", "0.005504993956671564", "0.005491302286152889", "0.005477644668686855", "0.005464021019578845", "0.00545043125434492", "0.0054368752887112345", "0.005423353038613559", "0.005409864420196741", "0.005396409349814191", "0.005382987744027348", "0.005369599519605185", "0.005356244593523682", "0.005342922882965306", "0.005329634305318512", "0.005316378778177204", "0.005303156219340258", "0.00528996654681099", "0.0052768096787966555", "0.00526368553370793", "0.005250594030158425", "0.005237535086964166", "0.0052245086231430945", "0.0052115145579145665", "0.005198552810698855", "0.005185623301116631", "0.005172725948988495", "0.005159860674334461", "0.005147027397373467", "0.005134226038522859", "0.00512145651839795", "0.005108718757811462", "0.005096012677773082", "0.00508333819948896", "0.005070695244361201", "0.0050580837339874105", "0.0050455035901601835", "0.00503295473486663", "0.005020437090287889", "0.005007950578798649", "0.004995495122966651", "0.004983070645552233", "0.004970677069507834", "0.004958314317977529", "0.004945982314296522", "0.004933680981990726", "0.004921410244776225", "0.004909170026558847", "0.0048969602514336765", "0.004884780843684585", "0.004872631727783748", "0.004860512828391204", "0.004848424070354368", "0.004836365378707559", "0.004824336678671571", "0.004812337895653155", "0.004800368955244605", "0.004788429783223271", "0.00477652030555111", "0.004764640448374205", "0.004752790138022353", "0.004740969301008549", "0.004729177864028579", "0.00471741575396054", "0.004705682897864399", "0.004693979222981524", "0.004682304656734251", "0.004670659126725434", "0.004659042560737964", "0.004647454886734382", "0.004635896032856363", "0.004624365927424321", "0.004612864498936943", "0.004601391676070756", "0.004589947387679656", "0.004578531562794525", "0.004567144130622721", "0.004555785020547693", "0.0045444541621285145", "0.004533151485099465", "0.004521876919369567", "0.004510630395022186", "0.004499411842314571", "0.004488221191677435", "0.004477058373714522", "0.004465923319202159", "0.004454815959088859", "0.0044437362244948665", "0.004432684046711748", "0.004421659357201942", "0.0044106620875983635", "0.004399692169703959", "0.004388749535491295", "0.004377834117102127", "0.004366945846846989", "0.004356084657204758", "0.004345250480822254", "0.004334443250513811", "0.004323662899260869", "0.004312909360211533", "0.004302182566680207", "0.0042914824521471245", "0.004280808950257977", "0.004270161994823491", "0.004259541519818998", "0.004248947459384061", "0.004238379747822035", "0.004227838319599677", "0.004217323109346733", "0.0042068340518555385", "0.004196371082080595", "0.004185934135138193", "0.004175523146305997", "0.0041651380510226476", "0.0041547787848873405", "0.0041444452836594745", "0.004134137483258197", "0.004123855319762044", "0.004113598729408536", "0.0041033676485937795", "0.00409316201387206", "0.004082981761955475", "0.004072826829713528", "0.004062697154172719", "0.004052592672516201", "0.004042513322083334", "0.004032459040369336", "0.004022429765024883", "0.004012425433855724", "0.004002445984822279", "0.0039924913560392935", "0.0039825614857754085", "0.003972656312452811", "0.0039627757746468345", "0.003952919811085593", "0.003943088360649578", "0.003933281362371305", "0.003923498755434923", "0.003913740479175826", "0.003904006473080314", "0.003894296676785166", "0.0038846110300773075", "0.0038749494728934205", "0.0038653119453195706", "0.0038556983875908417", "0.003846108740090951", "0.0038365429433519", "0.003827000938053592", "0.003817482665023469", "0.003807988065236137", "0.003798517079813012", "0.0037890696500219455", "0.0037796457172768793", "0.0037702452231374336", "0.003760868109308611", "0.0037515143176403924", "0.0037421837901273646", "0.0037328764689084134", "0.003723592296266315", "0.0037143312146274035", "0.0037050931665611963", "0.003695878094780059", "0.0036866859421388356", "0.0036775166516345007", "0.0036683701664057948", "0.0036592464297328883", "0.0036501453850370158", "0.0036410669758801476", "0.003632011145964594", "0.0036229778391327033", "0.0036139669993665007", "0.0036049785707873284", "0.0035960124976555", "0.003587068724369972", "0.0035781471954679863", "0.00356924785562472", "0.0035603706496529605", "0.0035515155225027497", "0.0035426824192610483", "0.003533871285151386", "0.003525082065533537", "0.003516314705903171", "0.003507569151891519", "0.0034988453492650275", "0.003490143243925033", "0.003481462781907431", "0.003472803909382326", "0.0034641665726536986", "0.0034555507181590877", "0.003446956292469248", "0.0034383832422878215", "0.003429831514450996", "0.0034213010559271955", "0.0034127918138167398", "0.003404303735351509", "0.003395836767894633", "0.003387390858940155", "0.0033789659561127092", "0.0033705620071671867", "0.003362178959988425", "0.0033538167625908845", "0.003345475363118319", "0.0033371547098434364", "0.003328854751167626", "0.003320575435620593", "0.0033123167118600644", "0.0033040785286714523", "0.003295860834967555", "0.0032876635797882323", "0.0032794867123000808", "0.0032713301817961335", "0.0032631939376955373", "0.003255077929543243", "0.0032469821070096813", "0.0032389064198904676", "0.0032308508181060785", "0.0032228152517015563", "0.0032147996708461633", "0.0032068040258331227", "0.003198828267079274", "0.0031908723451247807", "0.003182936210632811", "0.0031750198143892508", "0.003167123107302383", "0.0031592460404025937", "0.003151388564842052", "0.003143550631894429", "0.003135732192954583", "0.0031279331995382525", "0.003120153603281772", "0.0031123933559417563", "0.003104652409394822", "0.003096930715637249", "0.0030892282267847336", "0.0030815448950720567", "0.0030738806728528006", "0.0030662355125990444", "0.003058609366901082", "0.003051002188467121", "0.0030434139301229904", "0.003035844544811842", "0.003028293985593872", "0.003020762205646019", "0.0030132491582616793", "0.003005754796850408", "0.0029982790749376416", "0.002990821946164416", "0.0029833833642870446", "0.0029759632831768703", "0.002968561656819967", "0.0029611784393168477", "0.002953813584882177", "0.0029464670478445017", "0.002939138782645958", "0.0029318287438419924", "0.002924536886101071", "0.0029172631642044138", "0.0029100075330457022", "0.002902769947630807", "0.002895550363077497", "0.002888348734615178", "0.0028811650175846045", "0.0028739991674375997", "0.0028668511397367856", "0.002859720890155316", "0.0028526083744765812", "0.0028455135485939433", "0.0028384363685104693", "0.0028313767903386505", "0.0028243347703001353", "0.002817310264725446", "0.0028103032300537253", "0.0028033136228324557", "0.0027963413997171946", "0.002789386517471294", "0.0027824489329656495", "0.0027755286031784206", "0.0027686254851947796", "0.0027617395362066087", "0.002754870713512285", "0.002748018974516383", "0.002741184276729403", "0.002734366577767545", "0.0027275658353524096", "0.002720782007310756", "0.002714015051574226", "0.0027072649261790987", "0.0027005315892660205", "0.0026938149990797487", "0.0026871151139688867", "0.002680431892385635", "0.0026737652928855277", "0.002667115274127186", "0.0026604817948720325", "0.0026538648139840704", "0.002647264290429615", "0.0026406801832770345", "0.0026341124516964945", "0.0026275610549597156", "0.0026210259524397177", "0.002614507103610557", "0.0026080044680470904", "0.0026015180054247155", "0.0025950476755191246", "0.0025885934382060475", "0.002582155253461015", "0.0025757330813591", "0.0025693268820746796", "0.002562936615881173", "0.002556562243150812", "0.0025502037243543903", "0.0025438610200610133", "0.002537534090937851", "0.002531222897749906", "0.0025249274013597646", "0.002518647562727346", "0.002512383342909673", "0.0025061347030606255", "0.0024999016044306988", "0.0024936840083667573", "0.002487481876311808", "0.0024812951698047524", "0.0024751238504801517", "0.0024689678800679815", "0.002462827220393403", "0.0024567018333765287", "0.002450591681032179", "0.0024444967254696353", "0.0024384169288924388", "0.0024323522535981226", "0.002426302661977997", "0.0024202681165169044", "0.0024142485797929974", "0.002408244014477502", "0.0024022543833344813", "0.0023962796492206125", "0.002390319775084955", "0.0023843747239687177", "0.002378444459005027", "0.002372528943418707", "0.0023666281405260443", "0.0023607420137345706", "0.00235487052654281", "0.00234901364254009", "0.0023431713254062868", "0.002337343538911613", "0.0023315302469163837", "0.0023257314133708056", "0.0023199470023147423", "0.0023141769778774984", "0.002308421304277588", "0.002302679945822523", "0.0022969528669085897", "0.002291240032020618", "0.002285541405731775", "0.0022798569527033357", "0.002274186637684478", "0.002268530425512031", "0.0022628882811103024", "0.0022572601694908255", "0.0022516460557521606", "0.0022460459050796648", "0.002240459682745292", "0.0022348873541073655", "0.0022293288846103702", "0.0022237842397847297", "0.0022182533852466023", "0.0022127362866976668", "0.0022072329099248967", "0.002201743220800368", "0.0021962671852810297", "0.002190804769408513", "0.002185355939308889", "0.002179920661192491", "0.0021744989013536926", "0.0021690906261706954", "0.002163695802105317", "0.002158314395702796", "0.0021529463735915767", "0.002147591702483103", "0.0021422503491716075", "0.002136922280533915", "0.002131607463529231", "0.002126305865198939", "0.002121017452666391", "0.0021157421931367114", "0.0021104800538965904", "0.0021052310023140764", "0.0020999950058383805", "0.0020947720319996754", "0.002089562048408888", "0.002084365022757497", "0.002079180922817343", "0.0020740097164404186", "0.0020688513715586775", "0.0020637058561838234", "0.0020585731384071258", "0.002053453186399213", "0.00204834596840988", "0.002043251452767883", "0.0020381696078807534", "0.002033100402234596", "0.0020280438043939015", "0.002022999783001329", "0.002017968306777544", "0.002012949344521004", "0.0020079428651077567", "0.0020029488374912765", "0.0019979672307022457", "0.0019929980138483757", "0.001988041156114204", "0.0019830966267609163", "0.0019781643951261503", "0.0019732444306238043", "0.0019683367027438442", "0.001963441181052124", "0.001958557835190187", "0.001953686634875093", "0.001948827549899202", "0.0019439805501300148", "0.0019391456055099822", "0.0019343226860562947", "0.001929511761860731", "0.0019247128030894472", "0.0019199257799828032", "0.0019151506628551714", "0.00191038742209476", "0.0019056360281634245", "0.0019008964515964883", "0.0018961686630025515", "0.0018914526330633195", "0.0018867483325334157", "0.0018820557322402017", "0.00187737480308359", "0.0018727055160358732", "0.0018680478421415428", "0.0018634017525171029", "0.001858767218350892", "0.0018541442109029117", "0.001849532701504644", "0.0018449326615588685", "0.0018403440625394953", "0.0018357668759913805", "0.001831201073530154", "0.0018266466268420363", "0.0018221035076836736", "0.001817571687881955", "0.001813051139333842", "0.001808541834006187", "0.0018040437439355676", "0.0017995568412281146", "0.001795081098059332", "0.0017906164866739176", "0.0017861629793856156", "0.0017817205485770205", "0.0017772891666994195", "0.0017728688062726113", "0.0017684594398847473", "0.001764061040192155", "0.0017596735799191659", "0.001755297031857953", "0.0017509313688683584", "0.0017465765638777267", "0.001742232589880731", "0.0017378994199392156", "0.0017335770271820195", "0.0017292653848048228", "0.0017249644660699555", "0.0017206742443062635", "0.0017163946929089197", "0.0017121257853392698", "0.0017078674951246605", "0.001703619795858284", "0.0016993826611990095", "0.0016951560648712164", "0.0016909399806646387", "0.0016867343824341983", "0.0016825392440998445", "0.0016783545396463868", "0.0016741802431233428", "0.0016700163286447686", "0.001665862770389111", "0.0016617195425990224", "0.001657586619581233", "0.0016534639757063677", "0.0016493515854087985", "0.0016452494231864775", "0.001641157463600789", "0.001637075681276385", "0.0016330040509010303", "0.0016289425472254414", "0.001624891145063137", "0.001620849819290277", "0.0016168185448455056", "0.0016127972967298003", "0.0016087860500063127", "0.0016047847798002226", "0.0016007934612985643", "0.0015968120697500937", "0.0015928405804651279", "0.0015888789688153875", "0.0015849272102338443", "0.001580985280214576", "0.0015770531543126084", "0.0015731308081437668", "0.001569218217384519", "0.0015653153577718328", "0.00156142220510302", "0.0015575387352355897", "0.0015536649240870917", "0.0015498007476349772", "0.001545946181916444", "0.0015421012030282847", "0.0015382657871267455", "0.0015344399104273779", "0.0015306235492048854", "0.0015268166797929776", "0.0015230192785842286", "0.0015192313220299266", "0.00151545278663993", "0.0015116836489825162", "0.0015079238856842443", "0.0015041734734298055", "0.0015004323889618802", "0.0014967006090809893", "0.0014929781106453575", "0.0014892648705707666", "0.0014855608658304084", "0.0014818660734547471", "0.001478180470531379", "0.0014745040342048848", "0.0014708367416766818", "0.0014671785702049026", "0.001463529497104235", "0.001459889499745791", "0.0014562585555569602", "0.001452636642021277", "0.001449023736678276", "0.0014454198171233547", "0.0014418248610076313", "0.0014382388460378117", "0.0014346617499760462", "0.0014310935506397992", "0.0014275342259016956", "0.0014239837536894014", "0.0014204421119854828", "0.0014169092788272547", "0.001413385232306668", "0.0014098699505701556", "0.001406363411818506", "0.0014028655943067222", "0.0013993764763438924", "0.0013958960362930528", "0.001392424252571054", "0.0013889611036484245", "0.0013855065680492419", "0.0013820606243509967", "0.0013786232511844613", "0.001375194427233553", "0.0013717741312352066", "0.001368362341979244", "0.0013649590383082379", "0.0013615641991173786", "0.0013581778033543517", "0.0013547998300192025", "0.0013514302581642023", "0.0013480690668937255", "0.0013447162353641166", "0.0013413717427835613", "0.0013380355684119542", "0.0013347076915607773", "0.0013313880915929656", "0.0013280767479227835", "0.0013247736400156908", "0.0013214787473882221", "0.0013181920496078596", "0.0013149135262929023", "0.001311643157112335", "0.0013083809217857181", "0.0013051268000830484", "0.0013018807718246344", "0.0012986428168809787", "0.0012954129151726468", "0.0012921910466701457", "0.0012889771913937949", "0.0012857713294136101", "0.001282573440849174", "0.001279383505869516", "0.0012762015046929843", "0.00127302741758713", "0.0012698612248685797", "0.00126670290690292", "0.0012635524441045605", "0.001260409816936634", "0.0012572750059108581", "0.0012541479915874234", "0.0012510287545748659", "0.001247917275529954", "0.001244813535157566", "0.0012417175142105665", "0.0012386291934896932", "0.001235548553843434", "0.00123247557616791", "0.0012294102414067542", "0.001226352530550997", "0.0012233024246389459", "0.0012202599047560735", "0.0012172249520348841", "0.0012141975476548201", "0.001211177672842127", "0.0012081653088697446", "0.001205160437057188", "0.0012021630387704352", "0.0011991730954218087", "0.0011961905884698622", "0.0011932154994192614", "0.0011902478098206753", "0.0011872875012706595", "0.001184334555411538", "0.0011813889539312957", "0.00117845067856346", "0.0011755197110869951", "0.0011725960333261727", "0.0011696796271504805", "0.001166770474474494", "0.0011638685572577712", "0.0011609738575047374", "0.001158086357264577", "0.0011552060386311204", "0.0011523328837427338", "0.0011494668747822042", "0.0011466079939766362", "0.001143756223597338", "0.0011409115459597079", "0.0011380739434231314", "0.0011352433983908671", "0.0011324198933099438", "0.0011296034106710372", "0.0011267939330083783", "0.0011239914428996384", "0.0011211959229658179", "0.00111840735587114", "0.0011156257243229468", "0.0011128510110715887", "0.0011100831989103198", "0.001107322270675186", "0.0011045682092449256", "0.001101820997540859", "0.0010990806185267844", "0.0010963470552088684", "0.0010936202906355465", "0.001090900307897415", "0.0010881870901271234", "0.0010854806204992746", "0.0010827808822303207", "0.0010800878585784542", "0.0010774015328435052", "0.0010747218883668424", "0.0010720489085312653", "0.0010693825767609045", "0.0010667228765211133", "0.0010640697913183723", "0.0010614233047001828", "0.001058783400254966", "0.0010561500616119593", "0.0010535232724411178", "0.001050903016453011", "0.0010482892773987264", "0.0010456820390697555", "0.0010430812852979124", "0.0010404869999552202", "0.0010378991669538094", "0.001035317770245831", "0.0010327427938233455", "0.0010301742217182284", "0.0010276120380020677", "0.0010250562267860696", "0.0010225067722209583", "0.0010199636584968766", "0.0010174268698432876", "0.0010148963905288791", "0.0010123722048614638", "0.0010098542971878873", "0.0010073426518939187", "0.001004837253404167", "0.0010023380861819819", "0.000999845134729347", "0.000997358383586799", "0.000994877817333321", "0.0009924034205862516", "0.0009899351780011854", "0.0009874730742718838", "0.0009850170941301751", "0.0009825672223458639", "0.0009801234437266304", "0.0009776857431179438", "0.0009752541054029627", "0.0009728285155024452", "0.0009704089583746509", "0.0009679954190152511", "0.0009655878824572377", "0.0009631863337708251", "0.0009607907580633588", "0.0009584011404792269", "0.0009560174661997652", "0.0009536397204431631", "0.0009512678884643769", "0.0009489019555550353", "0.0009465419070433491", "0.0009441877282940176", "0.0009418394047081426", "0.0009394969217231342", "0.000937160264812623", "0.0009348294194863657", "0.0009325043712901601", "0.0009301851058057553", "0.0009278716086507594", "0.0009255638654785468", "0.0009232618619781814", "0.0009209655838743159", "0.0009186750169271098", "0.0009163901469321362", "0.000914110959720299", "0.000911837441157743", "0.000909569577145763", "0.0009073073536207216", "0.0009050507565539589", "0.0009027997719517073", "0.0009005543858550005", "0.0008983145843395932", "0.0008960803535158694", "0.0008938516795287629", "0.0008916285485576585", "0.0008894109468163234", "0.0008871988605528083", "0.000884992276049369", "0.0008827911796223766", "0.0008805955576222375", "0.000878405396433307", "0.0008762206824738015", "0.0008740414021957196", "0.0008718675420847549", "0.0008696990886602139", "0.0008675360284749287", "0.0008653783481151789", "0.0008632260342006045", "0.0008610790733841276", "0.000858937452351859", "0.0008568011578230308", "0.0008546701765499018", "0.0008525444953176817", "0.0008504241009444447", "0.0008483089802810527", "0.0008461991202110703", "0.0008440945076506856", "0.0008419951295486251", "0.0008399009728860782", "0.0008378120246766141", "0.0008357282719660983", "0.0008336497018326175", "0.0008315763013863953", "0.0008295080577697179", "0.0008274449581568436", "0.0008253869897539343", "0.0008233341397989731", "0.0008212863955616818", "0.0008192437443434435", "0.0008172061734772263", "0.0008151736703275019", "0.0008131462222901696", "0.0008111238167924742", "0.000809106441292933", "0.0008070940832812549", "0.0008050867302782645", "0.0008030843698358213", "0.0008010869895367475", "0.0007990945769947484", "0.0007971071198543334", "0.0007951246057907435", "0.0007931470225098742", "0.0007911743577481967", "0.0007892065992726818", "0.0007872437348807277", "0.0007852857524000816", "0.0007833326396887654", "0.0007813843846349972", "0.0007794409751571216", "0.0007775023992035306", "0.0007755686447525912", "0.0007736396998125676", "0.0007717155524215513", "0.0007697961906473848", "0.000767881602587585", "0.0007659717763692735", "0.0007640667001491032", "0.0007621663621131816", "0.0007602707504769951", "0.0007583798534853463", "0.0007564936594122707", "0.0007546121565609694", "0.000752735333263733", "0.0007508631778818736", "0.000748995678805649", "0.0007471328244541932", "0.0007452746032754412", "0.0007434210037460617", "0.0007415720143713818", "0.0007397276236853212", "0.000737887820250311", "0.0007360525926572334", "0.000734221929525348", "0.0007323958195022141", "0.000730574251263632", "0.0007287572135135638", "0.0007269446949840677", "0.0007251366844352247", "0.000723333170655073", "0.000721534142459536", "0.000719739588692354", "0.0007179494982250125", "0.0007161638599566769", "0.0007143826628141215", "0.0007126058957516616", "0.0007108335477510829", "0.0007090656078215762", "0.000707302064999669", "0.0007055429083491555", "0.0007037881269610281", "0.0007020377099534135", "0.0007002916464715031", "0.0006985499256874838", "0.0006968125368004746", "0.0006950794690364571", "0.00069335071164821", "0.00069162625391524", "0.0006899060851437189", "0.000688190194666415", "0.000686478571842628", "0.0006847712060581206", "0.0006830680867250557", "0.0006813692032819312", "0.0006796745451935118", "0.0006779841019507614", "0.0006762978630707868", "0.0006746158180967644", "0.0006729379565978776", "0.0006712642681692538", "0.0006695947424318983", "0.0006679293690326313", "0.0006662681376440209", "0.0006646110379643223", "0.0006629580597174121", "0.0006613091926527261", "0.0006596644265451924", "0.000658023751195172", "0.000656387156428393", "0.0006547546320958908", "0.0006531261680739369", "0.0006515017542639881", "0.0006498813805926142", "0.0006482650370114407", "0.0006466527134970823", "0.0006450444000510859", "0.0006434400866998653", "0.0006418397634946382", "0.0006402434205113683", "0.000638651047850701", "0.0006370626356379034", "0.0006354781740228006", "0.0006338976531797182", "0.0006323210633074185", "0.0006307483946290434", "0.0006291796373920459", "0.0006276147818681403", "0.0006260538183532337", "0.0006244967371673698", "0.0006229435286546658", "0.0006213941831832563", "0.0006198486911452311", "0.0006183070429565765", "0.0006167692290571141", "0.0006152352399104446", "0.0006137050660038869", "0.000612178697848418", "0.0006106561259786161", "0.0006091373409526013", "0.0006076223333519788", "0.000606111093781774", "0.0006046036128703823", "0.0006030998812695078", "0.0006015998896541044", "0.000600103628722317", "0.0005986110891954277", "0.0005971222618177952", "0.0005956371373567988", "0.000594155706602779", "0.0005926779603689835", "0.0005912038894915089", "0.0005897334848292419", "0.000588266737263806", "0.000586803637699503", "0.0005853441770632573", "0.0005838883463045577", "0.000582436136395404", "0.0005809875383302506", "0.0005795425431259495", "0.0005781011418216935", "0.0005766633254789636", "0.0005752290851814719", "0.0005737984120351071", "0.000572371297167877", "0.0005709477317298568", "0.0005695277068931323", "0.0005681112138517457", "0.0005666982438216399", "0.0005652887880406059", "0.0005638828377682278", "0.0005624803842858267", "0.0005610814188964092", "0.0005596859329246137", "0.0005582939177166547", "0.000556905364640267", "0.0005555202650846593", "0.0005541386104604545", "0.0005527603921996387", "0.0005513856017555068", "0.0005500142306026121", "0.0005486462702367112", "0.0005472817121747123", "0.000545920547954621", "0.0005445627691354901", "0.0005432083672973656", "0.0005418573340412372", "0.0005405096609889801", "0.0005391653397833095", "0.0005378243620877282", "0.0005364867195864678", "0.0005351524039844472", "0.0005338214070072143", "0.000532493720400897", "0.0005311693359321511", "0.0005298482453881103", "0.0005285304405763352", "0.0005272159133247621", "0.0005259046554816512", "0.0005245966589155381", "0.0005232919155151827", "0.0005219904171895188", "0.0005206921558676021", "0.0005193971234985632", "0.0005181053120515579", "0.0005168167135157115", "0.0005155313199000774", "0.0005142491232335822", "0.0005129701155649778", "0.0005116942889627907", "0.0005104216355152759", "0.0005091521473303648", "0.0005078858165356187", "0.0005066226352781766", "0.0005053625957247105", "0.0005041056900613743", "0.0005028519104937567", "0.0005016012492468304", "0.0005003536985649068", "0.0004991092507115877", "0.0004978678979697159", "0.0004966296326413248", "0.0004953944470475983", "0.0004941623335288165", "0.0004929332844443092", "0.0004917072921724111", "0.0004904843491104126", "0.0004892644476745133", "0.0004880475802997739", "0.00048683373944007096", "0.00048562291756804905", "0.0004844151071750748", "0.0004832103007711883", "0.00048200849088505973", "0.0004808096700639406", "0.0004796138308736203", "0.00047842096589837416", "0.0004772310677409256", "0.00047604412902239423", "0.0004748601423822513", "0.0004736791004782758", "0.00047250099598650756", "0.0004713258216012023", "0.00047015357003478517", "0.0004689842340178075", "0.00046781780629890035", "0.00046665427964473044", "0.00046549364683995354", "0.00046433590068717205", "0.0004631810340068887", "0.00046202903963746435", "0.000460879910435068", "0.0004597336392736403", "0.0004585902190448434", "0.0004574496426580196", "0.0004563119030401454", "0.0004551769931357902", "0.00045404490590707117", "0.00045291563433360834", "0.00045178917141248384", "0.0004506655101581963", "0.00044954464360261875", "0.0004484265647949539", "0.000447311266801693", "0.00044619874270657113", "0.00044508898561052717", "0.00044398198863165525", "0.00044287774490516803", "0.00044177624758335237", "0.0004406774898355255", "0.00043958146484799265", "0.0004384881658240068", "0.0004373975859837252", "0.0004363097185641675", "0.0004352245568191729", "0.00043414209401936043", "0.0004330623234520858", "0.00043198523842139896", "0.0004309108322480047", "0.00042983909826921986", "0.00042877002983893246", "0.00042770362032755927", "0.0004266398631220066", "0.0004255787516256291", "0.0004245202792581873", "0.00042346443945580705", "0.0004224112256709406", "0.00042136063137232445", "0.0004203126500449396", "0.00041926727518996963", "0.00041822450032476266", "0.0004171843189827903", "0.00041614672471360575", "0.0004151117110828069", "0.00041407927167199423", "0.00041304940007873205", "0.0004120220899165074", "0.0004109973348146922", "0.0004099751284185035", "0.00040895546438896355", "0.00040793833640285793", "0.00040692373815270243", "0.0004059116633466986", "0.0004049021057086971", "0.00040389505897815746", "0.0004028905169101107", "0.00040188847327511987", "0.0004008889218592418", "0.000399891856463987", "0.00039889727090628373", "0.00039790515901843833", "0.00039691551464809597", "0.00039592833165820457", "0.0003949436039269751", "0.000393961325347846", "0.00039298148982944", "0.00039200409129553347", "0.00039102912368501344", "0.00039005658095184247", "0.0003890864570650192", "0.0003881187460085436", "0.00038715344178137754", "0.00038619053839740886", "0.00038523002988541253", "0.0003842719102890158", "0.0003833161736666601", "0.00038236281409156426", "0.0003814118256516873", "0.0003804632024496925", "0.0003795169386029123", "0.0003785730282433066", "0.0003776314655174334", "0.00037669224458640715", "0.00037575535962586524", "0.00037482080482593", "0.00037388857439117466", "0.00037295866254058625", "0.0003720310635075301", "0.00037110577153971324", "0.0003701827808991501", "0.0003692620858621262", "0.00036834368071916293", "0.0003674275597749809", "0.00036651371734846644", "0.00036560214777263677", "0.00036469284539460085", "0.00036378580457552907", "0.0003628810196906165", "0.00036197848512904755", "0.00036107819529396056", "0.00036018014460241515", "0.0003592843274853561", "0.0003583907383875795", "0.000357499371767697", "0.0003566102220981035", "0.0003557232838649415", "0.0003548385515680673", "0.0003539560197210162", "0.0003530756828509697", "0.00035219753549872056", "0.0003513215722186408", "0.0003504477875786433", "0.0003495761761601545", "0.00034870673255807616", "0.0003478394513807529", "0.0003469743272499398", "0.00034611135480076816", "0.0003452505286817128", "0.00034439184355455747", "0.0003435352940943638", "0.00034268087498943685", "0.0003418285809412931", "0.00034097840666462605", "0.00034013034688727526", "0.00033928439635019255", "0.00033844054980741094", "0.0003375988020260081", "0.0003367591477860795", "0.00033592158188070186", "0.0003350860991159028", "0.0003342526943106274", "0.00033342136229670645", "0.0003325920979188266", "0.00033176489603449445", "0.0003309397515140068", "0.0003301166592404201", "0.000329295614109517", "0.00032847661102977405", "0.000327659644922331", "0.0003268447107209613", "0.000326031803372037", "0.0003252209178344992", "0.00032441204907982847", "0.0003236051920920098", "0.000322800341867506", "0.0003219974934152225", "0.00032119664175647835", "0.00032039778192497707", "0.0003196009089667721", "0.0003188060179402382", "0.00031801310391604175", "0.0003172221619771089", "0.00031643318721859433", "0.00031564617474785154", "0.00031486111968440447", "0.000314078017159914", "0.0003132968623181487", "0.00031251765031495743", "0.0003117403763182348", "0.0003109650355078954", "0.00031019162307584084", "0.00030942013422593086", "0.000308650564173955", "0.0003078829081476023", "0.00030711716138642796", "0.0003063533191418303", "0.0003055913766770181", "0.0003048313292669779", "0.00030407317219845127", "0.0003033169007699016", "0.0003025625102914848", "0.00030180999608502094", "0.000301059353483967", "0.00030031057783338404", "0.00029956366448991294", "0.0002988186088217414", "0.00029807540620857727", "0.0002973340520416207", "0.00029659454172353497", "0.00029585687066841464", "0.0002951210343017629", "0.00029438702806045995", "0.0002936548473927342", "0.0002929244877581347", "0.0002921959446275048", "0.0002914692134829511", "0.0002907442898178167", "0.00029002116913665494", "0.0002892998469551979", "0.0002885803188003326", "0.0002878625802100699", "0.0002871466267335181", "0.00028643245393085724", "0.0002857200573733079", "0.0002850094326431061", "0.0002843005753334761", "0.00028359348104860243", "0.00028288814540360183", "0.0002821845640244966", "0.0002814827325481894", "0.0002807826466224329", "0.0002800843019058045", "0.00027938769406768063", "0.0002786928187882068", "0.00027799967175827446", "0.0002773082486794909", "0.00027661854526415405", "0.0002759305572352276", "0.0002752442803263111", "0.00027455971028161554", "0.0002738768428559372", "0.00027319567381463116", "0.0002725161989335834", "0.00027183841399918595", "0.0002711623148083121", "0.0002704878971682869", "0.0002698151568968653", "0.00026914408982220227", "0.000268474691782829", "0.00026780695862762806", "0.0002671408862158053", "0.0002664764704168649", "0.0002658137071105858", "0.00026515259218699307", "0.0002644931215463338", "0.000263835291099053", "0.0002631790967657654", "0.0002625245344772333", "0.000261871600174338", "0.0002612202898080583", "0.0002605705993394415", "0.0002599225247395822", "0.0002592760619895941", "0.0002586312070805864", "0.00025798795601364026", "0.00025734630479978154", "0.0002567062494599569", "0.00025606778602501115", "0.0002554309105356593", "0.00025479561904246376", "0.00025416190760581107", "0.0002535297722958844", "0.0002528992091926425", "0.00025227021438579224", "0.0002516427839747676", "0.0002510169140687019", "0.0002503926007864077", "0.0002497698402563489", "0.00024914862861661854", "0.0002485289620149162", "0.00024791083660852134", "0.0002472942485642706", "0.00024667919405853554", "0.0002460656692771966", "0.00024545367041562007", "0.0002448431936786365", "0.0002442342352805136", "0.00024362679144493662", "0.0002430208584049815", "0.0002424164324030932", "0.000241813509691063", "0.00024121208653000463", "0.00024061215919032994", "0.0002400137239517268", "0.00023941677710313732", "0.00023882131494273222", "0.0002382273337778892", "0.00023763482992517122", "0.00023704379971030087", "0.00023645423946814072", "0.00023586614554266786", "0.0002352795142869524", "0.00023469434206313614", "0.0002341106252424074", "0.0002335283602049799", "0.0002329475433400711", "0.00023236817104587893", "0.00023179023972955872", "0.00023121374580720166", "0.00023063868570381385", "0.00023006505585329164", "0.0002294928526984008", "0.0002289220726907556", "0.00022835271229079405", "0.00022778476796775916", "0.00022721823619967416", "0.00022665311347332194", "0.00022608939628422403", "0.0002255270811366185", "0.00022496616454343546", "0.00022440664302628016", "0.00022384851311540923", "0.0002232917713497065", "0.00022273641427666648", "0.00022218243845237022", "0.00022162984044146337", "0.00022107861681713587", "0.00022052876416110172", "0.00021998027906357508", "0.00021943315812325236", "0.00021888739794728818", "0.00021834299515127576", "0.0002177999463592265", "0.0002172582482035487", "0.00021671789732502416", "0.00021617889037279164", "0.00021564122400432405", "0.00021510489488540523", "0.00021456989969011411", "0.00021403623510080118", "0.00021350389780806756", "0.00021297288451074537", "0.00021244319191587833", "0.00021191481673869857", "0.00021138775570260957", "0.00021086200553916288", "0.00021033756298803917", "0.0002098144247970291", "0.0002092925877220109", "0.00020877204852693136", "0.0002082528039837865", "0.00020773485087260092", "0.00020721818598140685", "0.00020670280610622524", "0.00020618870805104686", "0.0002056758886278102", "0.00020516434465638303", "0.0002046540729645435", "0.0002041450703879582", "0.00020363733377016513", "0.0002031308599625519", "0.0002026256458243371", "0.00020212168822255193", "0.00020161898403201864", "0.00020111753013533223", "0.00020061732342284186", "0.00020011836079263077", "0.00019962063915049635", "0.00019912415540993176", "0.0001986289064921078", "0.00019813488932585123", "0.0001976421008476287", "0.0001971505380015253", "0.00019666019773922647", "0.00019617107702000035", "0.0001956831728106767", "0.00019519648208562928", "0.00019471100182675793", "0.0001942267290234679", "0.00019374366067265227", "0.0001932617937786742", "0.00019278112535334613", "0.0001923016524159138", "0.00019182337199303518", "0.00019134628111876467", "0.00019087037683453213", "0.00019039565618912698", "0.0001899221162386778", "0.000189449754046635", "0.0001889785666837535", "0.00018850855122807267", "0.0001880397047648993", "0.00018757202438679028", "0.0001871055071935328", "0.0001866401502921272", "0.00018617595079677019", "0.0001857129058288345", "0.0001852510125168537", "0.00018479026799650178", "0.000184330669410578", "0.0001838722139089866", "0.0001834148986487217", "0.00018295872079384732", "0.00018250367751548093", "0.0001820497659917767", "0.00018159698340790626", "0.00018114532695604193", "0.0001806947938353406", "0.00018024538125192426", "0.00017979708641886356", "0.00017934990655616166", "0.00017890383889073463", "0.00017845888065639695", "0.00017801502909384187", "0.00017757228145062556", "0.00017713063498115038", "0.00017669008694664752", "0.00017625063461515912", "0.00017581227526152217", "0.00017537500616735232", "0.00017493882462102535", "0.00017450372791766127", "0.0001740697133591083", "0.00017363677825392424", "0.00017320491991736198", "0.00017277413567135089", "0.00017234442284448106", "0.00017191577877198765", "0.00017148820079573252", "0.00017106168626418867", "0.00017063623253242452", "0.00017021183696208666", "0.0001697884969213831", "0.00016936620978506747", "0.00016894497293442357", "0.00016852478375724753", "0.0001681056396478323", "0.00016768753800695251", "0.00016727047624184621", "0.0001668544517662012", "0.00016643946200013687", "0.0001660255043701892", "0.0001656125763092955", "0.00016520067525677696", "0.00016478979865832343", "0.00016437994396597828", "0.00016397110863812235", "0.000163563290139456", "0.00016315648594098702", "0.00016275069352001285", "0.00016234591036010462", "0.00016194213395109223", "0.00016153936178904955", "0.00016113759137627689", "0.0001607368202212878", "0.00016033704583879173", "0.0001599382657496793", "0.00015954047748100765", "0.00015914367856598462", "0.0001587478665439518", "0.0001583530389603723", "0.00015795919336681407", "0.00015756632732093296", "0.00015717443838646092", "0.00015678352413318896", "0.00015639358213695177", "0.00015600460997961335", "0.00015561660524905267", "0.0001552295655391469", "0.00015484348844975872", "0.00015445837158671938", "0.0001540742125618148", "0.0001536910089927715", "0.00015330875850324023", "0.0001529274587227821", "0.0001525471072868543", "0.00015216770183679496", "0.000151789240019808", "0.00015141171948894914", "0.0001510351379031119", "0.00015065949292701185", "0.00015028478223117256", "0.00014991100349191227", "0.00014953815439132734", "0.0001491662326172802", "0.00014879523586338312", "0.00014842516182898456", "0.00014805600821915594", "0.00014768777274467562", "0.00014732045312201554", "0.00014695404707332766", "0.0001465885523264292", "0.0001462239666147882", "0.00014586028767750973", "0.00014549751325932295", "0.00014513564111056523", "0.00014477466898716926", "0.00014441459465064986", "0.00014405541586808815", "0.00014369713041211983", "0.00014333973606091968", "0.0001429832305981884", "0.0001426276118131397", "0.00014227287750048507", "0.00014191902546042086", "0.00014156605349861537", "0.00014121395942619353", "0.0001408627410597252", "0.00014051239622120984", "0.0001401629227380649", "0.00013981431844311025", "0.0001394665811745569", "0.00013911970877599172", "0.00013877369909636494", "0.00013842854998997743", "0.00013808425931646602", "0.00013774082494079085", "0.00013739824473322303", "0.00013705651656932972", "0.00013671563832996195", "0.00013637560790124206", "0.0001360364231745489", "0.00013569808204650673", "0.00013536058241897026", "0.00013502392219901348", "0.00013468809929891484", "0.00013435311163614622", "0.0001340189571333582", "0.0001336856337183682", "0.000133353139324148", "0.00013302147188880972", "0.00013269062935559366", "0.00013236060967285627", "0.000132031410794056", "0.00013170303067774132", "0.00013137546728753883", "0.00013104871859213885", "0.00013072278256528482", "0.0001303976571857591", "0.000130073340437371", "0.00012974983030894494", "0.00012942712479430729", "0.0001291052218922737", "0.00012878411960663694", "0.0001284638159461554", "0.0001281443089245392", "0.00012782559656043864", "0.00012750767687743264", "0.00012719054790401505", "0.00012687420767358313", "0.00012655865422442594", "0.0001262438855997108", "0.0001259298998474728", "0.00012561669502060107", "0.00012530426917682766", "0.00012499262037871556", "0.00012468174669364655", "0.00012437164619380858", "0.0001240623169561844", "0.0001237537570625402", "0.00012344596459941236", "0.0001231389376580964", "0.00012283267433463562", "0.00012252717272980793", "0.00012222243094911565", "0.0001219184471027724", "0.00012161521930569189", "0.000121312745677477", "0.00012101102434240674", "0.00012071005342942529", "0.00012040983107213082", "0.00012011035540876375", "0.00011981162458219363", "0.00011951363673991026", "0.00011921639003401064", "0.00011891988262118735", "0.00011862411266271752", "0.00011832907832445205", "0.00011803477777680283", "0.00011774120919473294", "0.00011744837075774406", "0.00011715626064986561", "0.00011686487705964401", "0.00011657421818013124", "0.00011628428220887216", "0.00011599506734789578", "0.00011570657180370297", "0.000115418793787254", "0.00011513173151396", "0.00011484538320367034", "0.00011455974708066153", "0.00011427482137362653", "0.00011399060431566435", "0.00011370709414426775", "0.0001134242891013139", "0.00011314218743305201", "0.00011286078739009319", "0.00011258008722740005", "0.00011230008520427475", "0.00011202077958434883", "0.00011174216863557282", "0.00011146425063020524", "0.00011118702384480062", "0.00011091048656020106", "0.00011063463706152426", "0.0001103594736381527", "0.00011008499458372337", "0.00010981119819611783", "0.00010953808277745021", "0.00010926564663405836", "0.00010899388807649185", "0.00010872280541950219", "0.00010845239698203288", "0.00010818266108720791", "0.00010791359606232182", "0.00010764520023882983", "0.00010737747195233705", "0.00010711040954258776", "0.00010684401135345555", "0.00010657827573293359", "0.00010631320103312324", "0.00010604878561022439", "0.00010578502782452589", "0.00010552192604039398", "0.00010525947862626375", "0.00010499768395462758", "0.00010473654040202575", "0.00010447604634903683", "0.00010421620018026655", "0.00010395700028433838", "0.00010369844505388403", "0.00010344053288553221", "0.00010318326217990019", "0.00010292663134158238", "0.0001026706387791419", "0.00010241528290509928", "0.00010216056213592406", "0.00010190647489202366", "0.0001016530195977342", "0.0001014001946813112", "0.00010114799857491881", "0.00010089642971462057", "0.00010064548654037033", "0.0001003951674960014", "0.00010014547102921751", "9.989639559158371e-05", "9.964793963851548e-05", "9.940010162927062e-05", "9.915288002693825e-05", "9.890627329843071e-05", "9.866027991447263e-05", "9.841489834959287e-05", "9.817012708211378e-05", "9.792596459414239e-05", "9.768240937156141e-05", "9.743945990401885e-05", "9.719711468491922e-05", "9.695537221141459e-05", "9.671423098439433e-05", "9.647368950847631e-05", "9.623374629199814e-05", "9.59943998470067e-05", "9.575564868925029e-05", "9.551749133816822e-05", "9.52799263168822e-05", "9.504295215218745e-05", "9.480656737454325e-05", "9.457077051806351e-05", "9.433556012050796e-05", "9.410093472327367e-05", "9.386689287138491e-05", "9.363343311348472e-05", "9.340055400182631e-05", "9.316825409226318e-05", "9.293653194424059e-05", "9.270538612078716e-05", "9.24748151885048e-05", "9.224481771756114e-05", "9.201539228167948e-05", "9.178653745813048e-05", "9.155825182772367e-05", "9.133053397479826e-05", "9.110338248721411e-05", "9.087679595634325e-05", "9.065077297706164e-05", "9.04253121477395e-05", "9.020041207023308e-05", "8.997607134987651e-05", "8.975228859547199e-05", "8.952906241928245e-05", "8.930639143702184e-05", "8.908427426784703e-05", "8.886270953434968e-05", "8.864169586254683e-05", "8.842123188187275e-05", "8.820131622517084e-05", "8.798194752868477e-05", "8.77631244320498e-05", "8.754484557828454e-05", "8.732710961378314e-05", "8.710991518830579e-05", "8.689326095497101e-05", "8.667714557024758e-05", "8.646156769394526e-05", "8.624652598920765e-05", "8.603201912250282e-05", "8.581804576361552e-05", "8.560460458563938e-05", "8.539169426496779e-05", "8.517931348128614e-05", "8.496746091756387e-05", "8.475613526004626e-05", "8.454533519824515e-05", "8.433505942493262e-05", "8.412530663613193e-05", "8.391607553110912e-05", "8.370736481236539e-05", "8.349917318562943e-05", "8.329149935984834e-05", "8.308434204718088e-05", "8.287769996298837e-05", "8.267157182582722e-05", "8.246595635744123e-05", "8.22608522827536e-05", "8.205625832985787e-05", "8.185217323001193e-05", "8.164859571762917e-05", "8.144552453026978e-05", "8.12429584086347e-05", "8.104089609655679e-05", "8.083933634099283e-05", "8.063827789201616e-05", "8.043771950280922e-05", "8.023765992965492e-05", "8.003809793193002e-05", "7.983903227209647e-05", "7.964046171569414e-05", "7.944238503133356e-05", "7.924480099068753e-05", "7.904770836848383e-05", "7.885110594249795e-05", "7.86549924935452e-05", "7.845936680547292e-05", "7.826422766515316e-05", "7.806957386247563e-05", "7.787540419033932e-05", "7.76817174446454e-05", "7.748851242429031e-05", "7.729578793115717e-05", "7.710354277010953e-05", "7.691177574898303e-05", "7.672048567857839e-05", "7.652967137265442e-05", "7.633933164791985e-05", "7.614946532402644e-05", "7.59600712235619e-05", "7.577114817204235e-05", "7.558269499790468e-05", "7.539471053249969e-05", "7.520719361008512e-05", "7.502014306781768e-05", "7.483355774574627e-05", "7.464743648680508e-05", "7.446177813680559e-05", "7.427658154443043e-05", "7.409184556122532e-05", "7.390756904159231e-05", "7.372375084278316e-05", "7.354038982489135e-05", "7.33574848508455e-05", "7.317503478640266e-05", "7.299303850014037e-05", "7.28114948634507e-05", "7.263040275053221e-05", "7.244976103838399e-05", "7.226956860679767e-05", "7.208982433835149e-05", "7.191052711840251e-05", "7.173167583508007e-05", "7.155326937927923e-05", "7.137530664465318e-05", "7.119778652760675e-05", "7.102070792728993e-05", "7.084406974559031e-05", "7.066787088712663e-05", "7.049211025924237e-05", "7.031678677199809e-05", "7.014189933816568e-05", "6.99674468732206e-05", "6.979342829533621e-05", "6.961984252537598e-05", "6.944668848688785e-05", "6.927396510609668e-05", "6.910167131189796e-05", "6.892980603585151e-05", "6.875836821217415e-05", "6.858735677773345e-05", "6.841677067204151e-05", "6.824660883724761e-05", "6.80768702181321e-05", "6.790755376210011e-05", "6.773865841917428e-05", "6.757018314198916e-05", "6.740212688578385e-05", "6.723448860839594e-05", "6.706726727025528e-05", "6.690046183437722e-05", "6.673407126635603e-05", "6.656809453435868e-05", "6.64025306091188e-05", "6.62373784639296e-05", "6.607263707463784e-05", "6.590830541963784e-05", "6.574438247986447e-05", "6.558086723878711e-05", "6.541775868240377e-05", "6.525505579923394e-05", "6.509275758031328e-05", "6.493086301918653e-05", "6.476937111190159e-05", "6.460828085700362e-05", "6.444759125552847e-05", "6.428730131099635e-05", "6.412741002940587e-05", "6.396791641922817e-05", "6.380881949140011e-05", "6.365011825931852e-05", "6.349181173883436e-05", "6.333389894824585e-05", "6.31763789082933e-05", "6.301925064215222e-05", "6.286251317542763e-05", "6.270616553614835e-05", "6.255020675476025e-05", "6.239463586412065e-05", "6.223945189949249e-05", "6.208465389853825e-05", "6.193024090131323e-05", "6.177621195026089e-05", "6.162256609020617e-05", "6.14693023683494e-05", "6.131641983426072e-05", "6.116391753987436e-05", "6.1011794539482183e-05", "6.086004988972851e-05", "6.070868264960362e-05", "6.0557691880438226e-05", "6.040707664589783e-05", "6.025683601197684e-05", "6.010696904699205e-05", "5.9957474821578054e-05", "5.980835240868097e-05", "5.965960088355196e-05", "5.951121932374279e-05", "5.936320680909939e-05", "5.921556242175601e-05", "5.906828524612979e-05", "5.892137436891532e-05", "5.8774828879078326e-05", "5.862864786785079e-05", "5.848283042872463e-05", "5.8337375657446374e-05", "5.8192282652011844e-05", "5.804755051265997e-05", "5.79031783418675e-05", "5.775916524434369e-05", "5.761551032702456e-05", "5.74722126990667e-05", "5.732927147184299e-05", "5.718668575893631e-05", "5.704445467613399e-05", "5.690257734142252e-05", "5.676105287498238e-05", "5.661988039918188e-05", "5.647905903857252e-05", "5.633858791988285e-05", "5.619846617201338e-05", "5.605869292603145e-05", "5.591926731516527e-05", "5.578018847479881e-05", "5.564145554246667e-05", "5.5503067657848515e-05", "5.536502396276355e-05", "5.5227323601165393e-05", "5.508996571913705e-05", "5.4952949464885056e-05", "5.4816273988734456e-05", "5.467993844312386e-05", "5.4543941982599476e-05", "5.440828376381068e-05", "5.427296294550406e-05", "5.413797868851854e-05", "5.400333015578042e-05", "5.386901651229763e-05", "5.373503692515486e-05", "5.360139056350864e-05", "5.346807659858155e-05", "5.333509420365783e-05", "5.3202442554077494e-05", "5.307012082723197e-05", "5.293812820255826e-05", "5.2806463861534594e-05", "5.267512698767468e-05", "5.254411676652297e-05", "5.2413432385649814e-05", "5.2283073034645945e-05", "5.215303790511768e-05", "5.2023326190682185e-05", "5.1893937086961955e-05", "5.176486979158008e-05", "5.163612350415553e-05", "5.1507697426297574e-05", "5.1379590761601554e-05", "5.125180271564322e-05", "5.112433249597451e-05", "5.099717931211795e-05", "5.087034237556243e-05", "5.074382089975772e-05", "5.0617614100109834e-05", "5.049172119397646e-05", "5.0366141400661544e-05", "5.024087394141074e-05", "5.011591803940684e-05", "4.99912729197644e-05", "4.986693780952525e-05", "4.9742911937653897e-05", "4.9619194535032215e-05", "4.94957848344553e-05", "4.937268207062613e-05", "4.924988548015109e-05", "4.9127394301535405e-05", "4.900520777517822e-05", "4.8883325143367775e-05", "4.876174565027681e-05", "4.864046854195818e-05", "4.8519493066339644e-05", "4.8398818473219483e-05", "4.827844401426208e-05", "4.8158368942992777e-05", "4.803859251479349e-05", "4.791911398689837e-05", "4.7799932618388584e-05", "4.76810476701884e-05", "4.7562458405060015e-05", "4.744416408759925e-05", "4.732616398423112e-05", "4.720845736320517e-05", "4.709104349459072e-05", "4.6973921650272525e-05", "4.685709110394653e-05", "4.674055113111483e-05", "4.662430100908146e-05", "4.650834001694813e-05", "4.639266743560922e-05", "4.627728254774791e-05", "4.616218463783124e-05", "4.604737299210585e-05", "4.593284689859385e-05", "4.581860564708787e-05", "4.570464852914693e-05", "4.559097483809221e-05", "4.547758386900257e-05", "4.536447491870962e-05", "4.525164728579433e-05", "4.513910027058211e-05", "4.502683317513841e-05", "4.491484530326453e-05", "4.480313596049353e-05", "4.4691704454085434e-05", "4.458055009302347e-05", "4.446967218800931e-05", "4.4359070051459005e-05", "4.424874299749895e-05", "4.4138690341961164e-05", "4.402891140237929e-05", "4.391940549798451e-05", "4.381017194970126e-05", "4.3701210080142444e-05", "4.35925192136062e-05", "4.3484098676071145e-05", "4.3375947795192126e-05", "4.3268065900296206e-05", "4.316045232237874e-05", "4.305310639409866e-05", "4.294602744977499e-05", "4.283921482538217e-05", "4.273266785854614e-05", "4.2626385888540504e-05", "4.252036825628195e-05", "4.241461430432638e-05", "4.2309123376865024e-05", "4.2203894819720256e-05", "4.209892798034103e-05", "4.199422220779975e-05", "4.188977685278766e-05", "4.1785591267610814e-05", "4.168166480618613e-05", "4.1577996824037666e-05", "4.1474586678292084e-05", "4.137143372767524e-05", "4.126853733250774e-05", "4.116589685470111e-05", "4.1063511657754146e-05", "4.096138110674848e-05", "4.085950456834487e-05", "4.075788141077942e-05", "4.0656511003859525e-05", "4.0555392718959796e-05", "4.045452592901833e-05", "4.035391000853304e-05", "4.0253544333557296e-05", "4.0153428281696355e-05", "4.0053561232103635e-05", "3.9953942565476416e-05", "3.9854571664052536e-05", "3.97554479116061e-05", "3.9656570693443845e-05", "3.955793939640153e-05", "3.945955340883973e-05", "3.9361412120640285e-05", "3.926351492320264e-05", "3.916586120943967e-05", "3.906845037377442e-05", "3.897128181213582e-05", "3.8874354921955474e-05", "3.877766910216345e-05", "3.8681223753184774e-05", "3.858501827693588e-05", "3.848905207682046e-05", "3.8393324557726286e-05", "3.8297835126021054e-05", "3.820258318954892e-05", "3.810756815762698e-05", "3.801278944104126e-05", "3.7918246452043254e-05", "3.782393860434644e-05", "3.772986531312221e-05", "3.76360259949968e-05", "3.7542420068047066e-05", "3.744904695179748e-05", "3.735590606721595e-05", "3.7262996836710815e-05");
begin
    process(address)
    begin
        data_out <= to_stdlogicvector(lut(to_integer(unsigned(address))));
    end process;
end;

-- Add other necessary VHDL configurations and architectures if needed
